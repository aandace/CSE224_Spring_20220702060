magic
tech sky130A
magscale 1 2
timestamp 1745699999
<< nwell >>
rect 1066 2159 6662 7633
<< obsli1 >>
rect 1104 2159 6624 7633
<< obsm1 >>
rect 842 2128 6750 7664
<< metal2 >>
rect 2594 9077 2650 9877
rect 3238 9077 3294 9877
rect 3882 9077 3938 9877
rect 4526 9077 4582 9877
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
<< obsm2 >>
rect 846 9021 2538 9194
rect 2706 9021 3182 9194
rect 3350 9021 3826 9194
rect 3994 9021 4470 9194
rect 4638 9021 6744 9194
rect 846 856 6744 9021
rect 846 800 2538 856
rect 2706 800 3182 856
rect 3350 800 3826 856
rect 3994 800 4470 856
rect 4638 800 6744 856
<< metal3 >>
rect 0 7488 800 7608
rect 0 6808 800 6928
rect 0 6128 800 6248
rect 0 5448 800 5568
rect 6933 5448 7733 5568
rect 6933 4768 7733 4888
rect 6933 4088 7733 4208
rect 6933 3408 7733 3528
<< obsm3 >>
rect 880 7408 6938 7649
rect 798 7008 6938 7408
rect 880 6728 6938 7008
rect 798 6328 6938 6728
rect 880 6048 6938 6328
rect 798 5648 6938 6048
rect 880 5368 6853 5648
rect 798 4968 6938 5368
rect 798 4688 6853 4968
rect 798 4288 6938 4688
rect 798 4008 6853 4288
rect 798 3608 6938 4008
rect 798 3328 6853 3608
rect 798 2143 6938 3328
<< metal4 >>
rect 1633 2128 1953 7664
rect 2293 2128 2613 7752
rect 3012 2128 3332 7664
rect 3672 2128 3992 7752
rect 4391 2128 4711 7664
rect 5051 2128 5371 7752
rect 5770 2128 6090 7664
rect 6430 2128 6750 7752
<< obsm4 >>
rect 6867 5475 6933 5813
<< metal5 >>
rect 1056 7432 6750 7752
rect 1056 6772 6672 7092
rect 1056 6073 6750 6393
rect 1056 5413 6672 5733
rect 1056 4714 6750 5034
rect 1056 4054 6672 4374
rect 1056 3355 6750 3675
rect 1056 2695 6672 3015
<< labels >>
rlabel metal4 s 2293 2128 2613 7752 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 3672 2128 3992 7752 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 5051 2128 5371 7752 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 6430 2128 6750 7752 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 3355 6750 3675 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 4714 6750 5034 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 6073 6750 6393 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 7432 6750 7752 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 1633 2128 1953 7664 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 3012 2128 3332 7664 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 4391 2128 4711 7664 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 5770 2128 6090 7664 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 2695 6672 3015 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 4054 6672 4374 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 5413 6672 5733 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 6772 6672 7092 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 0 7488 800 7608 6 in[0]
port 3 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 in[1]
port 4 nsew signal input
rlabel metal2 s 2594 9077 2650 9877 6 in[2]
port 5 nsew signal input
rlabel metal2 s 3238 9077 3294 9877 6 in[3]
port 6 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 in[4]
port 7 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 in[5]
port 8 nsew signal input
rlabel metal3 s 6933 4088 7733 4208 6 in[6]
port 9 nsew signal input
rlabel metal3 s 6933 5448 7733 5568 6 in[7]
port 10 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 out[0]
port 11 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 out[1]
port 12 nsew signal output
rlabel metal2 s 4526 9077 4582 9877 6 out[2]
port 13 nsew signal output
rlabel metal2 s 3882 9077 3938 9877 6 out[3]
port 14 nsew signal output
rlabel metal2 s 2594 0 2650 800 6 out[4]
port 15 nsew signal output
rlabel metal2 s 3882 0 3938 800 6 out[5]
port 16 nsew signal output
rlabel metal3 s 6933 3408 7733 3528 6 out[6]
port 17 nsew signal output
rlabel metal3 s 6933 4768 7733 4888 6 out[7]
port 18 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 7733 9877
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 211792
string GDS_FILE /openlane/designs/twos_complement/runs/RUN_2025.04.26_20.39.24/results/signoff/twos_complement.magic.gds
string GDS_START 98260
<< end >>

