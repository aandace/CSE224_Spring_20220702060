magic
tech sky130A
magscale 1 2
timestamp 1745700003
<< checkpaint >>
rect -3932 -3932 11665 13809
<< viali >>
rect 4169 7497 4203 7531
rect 4813 7497 4847 7531
rect 1409 7361 1443 7395
rect 1685 7361 1719 7395
rect 2697 7361 2731 7395
rect 3341 7361 3375 7395
rect 4077 7361 4111 7395
rect 4721 7361 4755 7395
rect 1593 7157 1627 7191
rect 1869 7157 1903 7191
rect 2881 7157 2915 7191
rect 3525 7157 3559 7191
rect 4537 6953 4571 6987
rect 4353 6749 4387 6783
rect 2973 6409 3007 6443
rect 3801 6409 3835 6443
rect 3893 6409 3927 6443
rect 4629 6409 4663 6443
rect 3065 6341 3099 6375
rect 1869 6273 1903 6307
rect 2329 6273 2363 6307
rect 2605 6273 2639 6307
rect 2789 6273 2823 6307
rect 3341 6273 3375 6307
rect 3709 6273 3743 6307
rect 4261 6273 4295 6307
rect 4445 6273 4479 6307
rect 1777 6205 1811 6239
rect 3157 6205 3191 6239
rect 4169 6205 4203 6239
rect 1501 6069 1535 6103
rect 2145 6069 2179 6103
rect 2605 6069 2639 6103
rect 3065 6069 3099 6103
rect 3525 6069 3559 6103
rect 1501 5865 1535 5899
rect 2973 5865 3007 5899
rect 3065 5729 3099 5763
rect 1685 5661 1719 5695
rect 1777 5661 1811 5695
rect 2789 5661 2823 5695
rect 2881 5661 2915 5695
rect 6285 5661 6319 5695
rect 1961 5525 1995 5559
rect 6101 5525 6135 5559
rect 5273 5185 5307 5219
rect 5917 5185 5951 5219
rect 5181 5117 5215 5151
rect 5641 5117 5675 5151
rect 6101 4981 6135 5015
rect 6285 4573 6319 4607
rect 6101 4437 6135 4471
rect 2881 4097 2915 4131
rect 3065 4097 3099 4131
rect 2881 3893 2915 3927
rect 2789 3689 2823 3723
rect 4169 3621 4203 3655
rect 5181 3621 5215 3655
rect 5733 3621 5767 3655
rect 3157 3553 3191 3587
rect 5365 3553 5399 3587
rect 2513 3485 2547 3519
rect 2605 3485 2639 3519
rect 3065 3485 3099 3519
rect 3985 3485 4019 3519
rect 4077 3485 4111 3519
rect 4261 3485 4295 3519
rect 5549 3485 5583 3519
rect 6009 3485 6043 3519
rect 4445 3417 4479 3451
rect 4905 3417 4939 3451
rect 3433 3349 3467 3383
rect 6193 3349 6227 3383
rect 3065 3145 3099 3179
rect 4629 3145 4663 3179
rect 2973 3009 3007 3043
rect 3157 3009 3191 3043
rect 4169 3009 4203 3043
rect 4353 3009 4387 3043
rect 4445 3009 4479 3043
rect 4169 2805 4203 2839
rect 3525 2601 3559 2635
rect 4629 2601 4663 2635
rect 2973 2397 3007 2431
rect 3341 2397 3375 2431
rect 3985 2397 4019 2431
rect 4813 2397 4847 2431
rect 2789 2261 2823 2295
rect 4169 2261 4203 2295
<< metal1 >>
rect 1104 7642 6750 7664
rect 1104 7590 2299 7642
rect 2351 7590 2363 7642
rect 2415 7590 2427 7642
rect 2479 7590 2491 7642
rect 2543 7590 2555 7642
rect 2607 7590 3678 7642
rect 3730 7590 3742 7642
rect 3794 7590 3806 7642
rect 3858 7590 3870 7642
rect 3922 7590 3934 7642
rect 3986 7590 5057 7642
rect 5109 7590 5121 7642
rect 5173 7590 5185 7642
rect 5237 7590 5249 7642
rect 5301 7590 5313 7642
rect 5365 7590 6436 7642
rect 6488 7590 6500 7642
rect 6552 7590 6564 7642
rect 6616 7590 6628 7642
rect 6680 7590 6692 7642
rect 6744 7590 6750 7642
rect 1104 7568 6750 7590
rect 4062 7488 4068 7540
rect 4120 7528 4126 7540
rect 4157 7531 4215 7537
rect 4157 7528 4169 7531
rect 4120 7500 4169 7528
rect 4120 7488 4126 7500
rect 4157 7497 4169 7500
rect 4203 7497 4215 7531
rect 4157 7491 4215 7497
rect 4798 7488 4804 7540
rect 4856 7488 4862 7540
rect 842 7352 848 7404
rect 900 7392 906 7404
rect 1397 7395 1455 7401
rect 1397 7392 1409 7395
rect 900 7364 1409 7392
rect 900 7352 906 7364
rect 1397 7361 1409 7364
rect 1443 7361 1455 7395
rect 1397 7355 1455 7361
rect 1486 7352 1492 7404
rect 1544 7392 1550 7404
rect 1673 7395 1731 7401
rect 1673 7392 1685 7395
rect 1544 7364 1685 7392
rect 1544 7352 1550 7364
rect 1673 7361 1685 7364
rect 1719 7361 1731 7395
rect 1673 7355 1731 7361
rect 2682 7352 2688 7404
rect 2740 7352 2746 7404
rect 3326 7352 3332 7404
rect 3384 7352 3390 7404
rect 4062 7352 4068 7404
rect 4120 7352 4126 7404
rect 4709 7395 4767 7401
rect 4709 7361 4721 7395
rect 4755 7392 4767 7395
rect 4798 7392 4804 7404
rect 4755 7364 4804 7392
rect 4755 7361 4767 7364
rect 4709 7355 4767 7361
rect 4798 7352 4804 7364
rect 4856 7352 4862 7404
rect 1394 7148 1400 7200
rect 1452 7188 1458 7200
rect 1581 7191 1639 7197
rect 1581 7188 1593 7191
rect 1452 7160 1593 7188
rect 1452 7148 1458 7160
rect 1581 7157 1593 7160
rect 1627 7157 1639 7191
rect 1581 7151 1639 7157
rect 1857 7191 1915 7197
rect 1857 7157 1869 7191
rect 1903 7188 1915 7191
rect 2038 7188 2044 7200
rect 1903 7160 2044 7188
rect 1903 7157 1915 7160
rect 1857 7151 1915 7157
rect 2038 7148 2044 7160
rect 2096 7148 2102 7200
rect 2866 7148 2872 7200
rect 2924 7148 2930 7200
rect 3510 7148 3516 7200
rect 3568 7148 3574 7200
rect 1104 7098 6624 7120
rect 1104 7046 1639 7098
rect 1691 7046 1703 7098
rect 1755 7046 1767 7098
rect 1819 7046 1831 7098
rect 1883 7046 1895 7098
rect 1947 7046 3018 7098
rect 3070 7046 3082 7098
rect 3134 7046 3146 7098
rect 3198 7046 3210 7098
rect 3262 7046 3274 7098
rect 3326 7046 4397 7098
rect 4449 7046 4461 7098
rect 4513 7046 4525 7098
rect 4577 7046 4589 7098
rect 4641 7046 4653 7098
rect 4705 7046 5776 7098
rect 5828 7046 5840 7098
rect 5892 7046 5904 7098
rect 5956 7046 5968 7098
rect 6020 7046 6032 7098
rect 6084 7046 6624 7098
rect 1104 7024 6624 7046
rect 4525 6987 4583 6993
rect 4525 6953 4537 6987
rect 4571 6984 4583 6987
rect 4798 6984 4804 6996
rect 4571 6956 4804 6984
rect 4571 6953 4583 6956
rect 4525 6947 4583 6953
rect 4798 6944 4804 6956
rect 4856 6944 4862 6996
rect 4341 6783 4399 6789
rect 4341 6749 4353 6783
rect 4387 6780 4399 6783
rect 4614 6780 4620 6792
rect 4387 6752 4620 6780
rect 4387 6749 4399 6752
rect 4341 6743 4399 6749
rect 4614 6740 4620 6752
rect 4672 6740 4678 6792
rect 1104 6554 6750 6576
rect 1104 6502 2299 6554
rect 2351 6502 2363 6554
rect 2415 6502 2427 6554
rect 2479 6502 2491 6554
rect 2543 6502 2555 6554
rect 2607 6502 3678 6554
rect 3730 6502 3742 6554
rect 3794 6502 3806 6554
rect 3858 6502 3870 6554
rect 3922 6502 3934 6554
rect 3986 6502 5057 6554
rect 5109 6502 5121 6554
rect 5173 6502 5185 6554
rect 5237 6502 5249 6554
rect 5301 6502 5313 6554
rect 5365 6502 6436 6554
rect 6488 6502 6500 6554
rect 6552 6502 6564 6554
rect 6616 6502 6628 6554
rect 6680 6502 6692 6554
rect 6744 6502 6750 6554
rect 1104 6480 6750 6502
rect 2961 6443 3019 6449
rect 2961 6409 2973 6443
rect 3007 6440 3019 6443
rect 3007 6412 3280 6440
rect 3007 6409 3019 6412
rect 2961 6403 3019 6409
rect 2682 6372 2688 6384
rect 1780 6344 2360 6372
rect 1394 6196 1400 6248
rect 1452 6236 1458 6248
rect 1780 6245 1808 6344
rect 1857 6307 1915 6313
rect 1857 6273 1869 6307
rect 1903 6304 1915 6307
rect 2038 6304 2044 6316
rect 1903 6276 2044 6304
rect 1903 6273 1915 6276
rect 1857 6267 1915 6273
rect 2038 6264 2044 6276
rect 2096 6264 2102 6316
rect 2332 6313 2360 6344
rect 2608 6344 2688 6372
rect 2608 6313 2636 6344
rect 2682 6332 2688 6344
rect 2740 6372 2746 6384
rect 3053 6375 3111 6381
rect 3053 6372 3065 6375
rect 2740 6344 3065 6372
rect 2740 6332 2746 6344
rect 3053 6341 3065 6344
rect 3099 6341 3111 6375
rect 3053 6335 3111 6341
rect 2317 6307 2375 6313
rect 2317 6273 2329 6307
rect 2363 6304 2375 6307
rect 2593 6307 2651 6313
rect 2593 6304 2605 6307
rect 2363 6276 2605 6304
rect 2363 6273 2375 6276
rect 2317 6267 2375 6273
rect 2593 6273 2605 6276
rect 2639 6273 2651 6307
rect 2593 6267 2651 6273
rect 2777 6307 2835 6313
rect 2777 6273 2789 6307
rect 2823 6304 2835 6307
rect 2866 6304 2872 6316
rect 2823 6276 2872 6304
rect 2823 6273 2835 6276
rect 2777 6267 2835 6273
rect 2866 6264 2872 6276
rect 2924 6264 2930 6316
rect 1765 6239 1823 6245
rect 1765 6236 1777 6239
rect 1452 6208 1777 6236
rect 1452 6196 1458 6208
rect 1765 6205 1777 6208
rect 1811 6205 1823 6239
rect 1765 6199 1823 6205
rect 2056 6168 2084 6264
rect 3145 6239 3203 6245
rect 3145 6236 3157 6239
rect 2608 6208 3157 6236
rect 2608 6168 2636 6208
rect 3145 6205 3157 6208
rect 3191 6205 3203 6239
rect 3252 6236 3280 6412
rect 3510 6400 3516 6452
rect 3568 6440 3574 6452
rect 3789 6443 3847 6449
rect 3789 6440 3801 6443
rect 3568 6412 3801 6440
rect 3568 6400 3574 6412
rect 3789 6409 3801 6412
rect 3835 6409 3847 6443
rect 3789 6403 3847 6409
rect 3881 6443 3939 6449
rect 3881 6409 3893 6443
rect 3927 6440 3939 6443
rect 4062 6440 4068 6452
rect 3927 6412 4068 6440
rect 3927 6409 3939 6412
rect 3881 6403 3939 6409
rect 4062 6400 4068 6412
rect 4120 6400 4126 6452
rect 4614 6400 4620 6452
rect 4672 6400 4678 6452
rect 3329 6307 3387 6313
rect 3329 6273 3341 6307
rect 3375 6304 3387 6307
rect 3528 6304 3556 6400
rect 3375 6276 3556 6304
rect 3697 6307 3755 6313
rect 3375 6273 3387 6276
rect 3329 6267 3387 6273
rect 3697 6273 3709 6307
rect 3743 6304 3755 6307
rect 4249 6307 4307 6313
rect 4249 6304 4261 6307
rect 3743 6276 4261 6304
rect 3743 6273 3755 6276
rect 3697 6267 3755 6273
rect 4249 6273 4261 6276
rect 4295 6273 4307 6307
rect 4249 6267 4307 6273
rect 4433 6307 4491 6313
rect 4433 6273 4445 6307
rect 4479 6273 4491 6307
rect 4433 6267 4491 6273
rect 3712 6236 3740 6267
rect 3252 6208 3740 6236
rect 3145 6199 3203 6205
rect 4154 6196 4160 6248
rect 4212 6196 4218 6248
rect 2056 6140 2636 6168
rect 2608 6112 2636 6140
rect 2866 6128 2872 6180
rect 2924 6168 2930 6180
rect 2924 6140 3096 6168
rect 2924 6128 2930 6140
rect 1486 6060 1492 6112
rect 1544 6060 1550 6112
rect 2130 6060 2136 6112
rect 2188 6060 2194 6112
rect 2590 6060 2596 6112
rect 2648 6060 2654 6112
rect 3068 6109 3096 6140
rect 3418 6128 3424 6180
rect 3476 6168 3482 6180
rect 4448 6168 4476 6267
rect 3476 6140 4476 6168
rect 3476 6128 3482 6140
rect 3053 6103 3111 6109
rect 3053 6069 3065 6103
rect 3099 6069 3111 6103
rect 3053 6063 3111 6069
rect 3513 6103 3571 6109
rect 3513 6069 3525 6103
rect 3559 6100 3571 6103
rect 4154 6100 4160 6112
rect 3559 6072 4160 6100
rect 3559 6069 3571 6072
rect 3513 6063 3571 6069
rect 4154 6060 4160 6072
rect 4212 6060 4218 6112
rect 1104 6010 6624 6032
rect 1104 5958 1639 6010
rect 1691 5958 1703 6010
rect 1755 5958 1767 6010
rect 1819 5958 1831 6010
rect 1883 5958 1895 6010
rect 1947 5958 3018 6010
rect 3070 5958 3082 6010
rect 3134 5958 3146 6010
rect 3198 5958 3210 6010
rect 3262 5958 3274 6010
rect 3326 5958 4397 6010
rect 4449 5958 4461 6010
rect 4513 5958 4525 6010
rect 4577 5958 4589 6010
rect 4641 5958 4653 6010
rect 4705 5958 5776 6010
rect 5828 5958 5840 6010
rect 5892 5958 5904 6010
rect 5956 5958 5968 6010
rect 6020 5958 6032 6010
rect 6084 5958 6624 6010
rect 1104 5936 6624 5958
rect 1210 5856 1216 5908
rect 1268 5896 1274 5908
rect 1489 5899 1547 5905
rect 1489 5896 1501 5899
rect 1268 5868 1501 5896
rect 1268 5856 1274 5868
rect 1489 5865 1501 5868
rect 1535 5865 1547 5899
rect 1489 5859 1547 5865
rect 2961 5899 3019 5905
rect 2961 5865 2973 5899
rect 3007 5896 3019 5899
rect 3418 5896 3424 5908
rect 3007 5868 3424 5896
rect 3007 5865 3019 5868
rect 2961 5859 3019 5865
rect 3418 5856 3424 5868
rect 3476 5856 3482 5908
rect 2866 5788 2872 5840
rect 2924 5828 2930 5840
rect 2924 5800 3096 5828
rect 2924 5788 2930 5800
rect 1486 5720 1492 5772
rect 1544 5760 1550 5772
rect 3068 5769 3096 5800
rect 3053 5763 3111 5769
rect 1544 5732 1808 5760
rect 1544 5720 1550 5732
rect 1780 5701 1808 5732
rect 3053 5729 3065 5763
rect 3099 5729 3111 5763
rect 3053 5723 3111 5729
rect 1673 5695 1731 5701
rect 1673 5661 1685 5695
rect 1719 5661 1731 5695
rect 1673 5655 1731 5661
rect 1765 5695 1823 5701
rect 1765 5661 1777 5695
rect 1811 5661 1823 5695
rect 1765 5655 1823 5661
rect 1688 5624 1716 5655
rect 2590 5652 2596 5704
rect 2648 5692 2654 5704
rect 2777 5695 2835 5701
rect 2777 5692 2789 5695
rect 2648 5664 2789 5692
rect 2648 5652 2654 5664
rect 2777 5661 2789 5664
rect 2823 5661 2835 5695
rect 2777 5655 2835 5661
rect 2869 5695 2927 5701
rect 2869 5661 2881 5695
rect 2915 5661 2927 5695
rect 2869 5655 2927 5661
rect 2130 5624 2136 5636
rect 1688 5596 2136 5624
rect 2130 5584 2136 5596
rect 2188 5584 2194 5636
rect 2682 5584 2688 5636
rect 2740 5624 2746 5636
rect 2884 5624 2912 5655
rect 6270 5652 6276 5704
rect 6328 5652 6334 5704
rect 2740 5596 2912 5624
rect 2740 5584 2746 5596
rect 1946 5516 1952 5568
rect 2004 5516 2010 5568
rect 5442 5516 5448 5568
rect 5500 5556 5506 5568
rect 6089 5559 6147 5565
rect 6089 5556 6101 5559
rect 5500 5528 6101 5556
rect 5500 5516 5506 5528
rect 6089 5525 6101 5528
rect 6135 5525 6147 5559
rect 6089 5519 6147 5525
rect 1104 5466 6750 5488
rect 1104 5414 2299 5466
rect 2351 5414 2363 5466
rect 2415 5414 2427 5466
rect 2479 5414 2491 5466
rect 2543 5414 2555 5466
rect 2607 5414 3678 5466
rect 3730 5414 3742 5466
rect 3794 5414 3806 5466
rect 3858 5414 3870 5466
rect 3922 5414 3934 5466
rect 3986 5414 5057 5466
rect 5109 5414 5121 5466
rect 5173 5414 5185 5466
rect 5237 5414 5249 5466
rect 5301 5414 5313 5466
rect 5365 5414 6436 5466
rect 6488 5414 6500 5466
rect 6552 5414 6564 5466
rect 6616 5414 6628 5466
rect 6680 5414 6692 5466
rect 6744 5414 6750 5466
rect 1104 5392 6750 5414
rect 5261 5219 5319 5225
rect 5261 5185 5273 5219
rect 5307 5216 5319 5219
rect 5442 5216 5448 5228
rect 5307 5188 5448 5216
rect 5307 5185 5319 5188
rect 5261 5179 5319 5185
rect 5442 5176 5448 5188
rect 5500 5176 5506 5228
rect 5905 5219 5963 5225
rect 5905 5216 5917 5219
rect 5644 5188 5917 5216
rect 4982 5108 4988 5160
rect 5040 5148 5046 5160
rect 5644 5157 5672 5188
rect 5905 5185 5917 5188
rect 5951 5185 5963 5219
rect 5905 5179 5963 5185
rect 5169 5151 5227 5157
rect 5169 5148 5181 5151
rect 5040 5120 5181 5148
rect 5040 5108 5046 5120
rect 5169 5117 5181 5120
rect 5215 5117 5227 5151
rect 5169 5111 5227 5117
rect 5629 5151 5687 5157
rect 5629 5117 5641 5151
rect 5675 5117 5687 5151
rect 5629 5111 5687 5117
rect 6089 5015 6147 5021
rect 6089 4981 6101 5015
rect 6135 5012 6147 5015
rect 6178 5012 6184 5024
rect 6135 4984 6184 5012
rect 6135 4981 6147 4984
rect 6089 4975 6147 4981
rect 6178 4972 6184 4984
rect 6236 4972 6242 5024
rect 1104 4922 6624 4944
rect 1104 4870 1639 4922
rect 1691 4870 1703 4922
rect 1755 4870 1767 4922
rect 1819 4870 1831 4922
rect 1883 4870 1895 4922
rect 1947 4870 3018 4922
rect 3070 4870 3082 4922
rect 3134 4870 3146 4922
rect 3198 4870 3210 4922
rect 3262 4870 3274 4922
rect 3326 4870 4397 4922
rect 4449 4870 4461 4922
rect 4513 4870 4525 4922
rect 4577 4870 4589 4922
rect 4641 4870 4653 4922
rect 4705 4870 5776 4922
rect 5828 4870 5840 4922
rect 5892 4870 5904 4922
rect 5956 4870 5968 4922
rect 6020 4870 6032 4922
rect 6084 4870 6624 4922
rect 1104 4848 6624 4870
rect 6270 4564 6276 4616
rect 6328 4564 6334 4616
rect 4798 4428 4804 4480
rect 4856 4468 4862 4480
rect 6089 4471 6147 4477
rect 6089 4468 6101 4471
rect 4856 4440 6101 4468
rect 4856 4428 4862 4440
rect 6089 4437 6101 4440
rect 6135 4437 6147 4471
rect 6089 4431 6147 4437
rect 1104 4378 6750 4400
rect 1104 4326 2299 4378
rect 2351 4326 2363 4378
rect 2415 4326 2427 4378
rect 2479 4326 2491 4378
rect 2543 4326 2555 4378
rect 2607 4326 3678 4378
rect 3730 4326 3742 4378
rect 3794 4326 3806 4378
rect 3858 4326 3870 4378
rect 3922 4326 3934 4378
rect 3986 4326 5057 4378
rect 5109 4326 5121 4378
rect 5173 4326 5185 4378
rect 5237 4326 5249 4378
rect 5301 4326 5313 4378
rect 5365 4326 6436 4378
rect 6488 4326 6500 4378
rect 6552 4326 6564 4378
rect 6616 4326 6628 4378
rect 6680 4326 6692 4378
rect 6744 4326 6750 4378
rect 1104 4304 6750 4326
rect 2774 4088 2780 4140
rect 2832 4128 2838 4140
rect 2869 4131 2927 4137
rect 2869 4128 2881 4131
rect 2832 4100 2881 4128
rect 2832 4088 2838 4100
rect 2869 4097 2881 4100
rect 2915 4097 2927 4131
rect 2869 4091 2927 4097
rect 3053 4131 3111 4137
rect 3053 4097 3065 4131
rect 3099 4128 3111 4131
rect 3418 4128 3424 4140
rect 3099 4100 3424 4128
rect 3099 4097 3111 4100
rect 3053 4091 3111 4097
rect 3418 4088 3424 4100
rect 3476 4088 3482 4140
rect 2866 3884 2872 3936
rect 2924 3884 2930 3936
rect 1104 3834 6624 3856
rect 1104 3782 1639 3834
rect 1691 3782 1703 3834
rect 1755 3782 1767 3834
rect 1819 3782 1831 3834
rect 1883 3782 1895 3834
rect 1947 3782 3018 3834
rect 3070 3782 3082 3834
rect 3134 3782 3146 3834
rect 3198 3782 3210 3834
rect 3262 3782 3274 3834
rect 3326 3782 4397 3834
rect 4449 3782 4461 3834
rect 4513 3782 4525 3834
rect 4577 3782 4589 3834
rect 4641 3782 4653 3834
rect 4705 3782 5776 3834
rect 5828 3782 5840 3834
rect 5892 3782 5904 3834
rect 5956 3782 5968 3834
rect 6020 3782 6032 3834
rect 6084 3782 6624 3834
rect 1104 3760 6624 3782
rect 2774 3680 2780 3732
rect 2832 3680 2838 3732
rect 4246 3720 4252 3732
rect 2976 3692 4252 3720
rect 2976 3652 3004 3692
rect 4246 3680 4252 3692
rect 4304 3680 4310 3732
rect 4062 3652 4068 3664
rect 2608 3624 3004 3652
rect 3068 3624 4068 3652
rect 2608 3525 2636 3624
rect 3068 3525 3096 3624
rect 4062 3612 4068 3624
rect 4120 3652 4126 3664
rect 4157 3655 4215 3661
rect 4157 3652 4169 3655
rect 4120 3624 4169 3652
rect 4120 3612 4126 3624
rect 4157 3621 4169 3624
rect 4203 3621 4215 3655
rect 4157 3615 4215 3621
rect 4982 3612 4988 3664
rect 5040 3652 5046 3664
rect 5169 3655 5227 3661
rect 5169 3652 5181 3655
rect 5040 3624 5181 3652
rect 5040 3612 5046 3624
rect 5169 3621 5181 3624
rect 5215 3621 5227 3655
rect 5169 3615 5227 3621
rect 5721 3655 5779 3661
rect 5721 3621 5733 3655
rect 5767 3621 5779 3655
rect 5721 3615 5779 3621
rect 3142 3544 3148 3596
rect 3200 3584 3206 3596
rect 3418 3584 3424 3596
rect 3200 3556 3424 3584
rect 3200 3544 3206 3556
rect 3418 3544 3424 3556
rect 3476 3544 3482 3596
rect 4338 3584 4344 3596
rect 3988 3556 4344 3584
rect 3988 3525 4016 3556
rect 4338 3544 4344 3556
rect 4396 3584 4402 3596
rect 4798 3584 4804 3596
rect 4396 3556 4804 3584
rect 4396 3544 4402 3556
rect 4798 3544 4804 3556
rect 4856 3544 4862 3596
rect 5353 3587 5411 3593
rect 5353 3553 5365 3587
rect 5399 3584 5411 3587
rect 5399 3556 5580 3584
rect 5399 3553 5411 3556
rect 5353 3547 5411 3553
rect 2501 3519 2559 3525
rect 2501 3485 2513 3519
rect 2547 3485 2559 3519
rect 2501 3479 2559 3485
rect 2593 3519 2651 3525
rect 2593 3485 2605 3519
rect 2639 3485 2651 3519
rect 2593 3479 2651 3485
rect 3053 3519 3111 3525
rect 3053 3485 3065 3519
rect 3099 3485 3111 3519
rect 3053 3479 3111 3485
rect 3973 3519 4031 3525
rect 3973 3485 3985 3519
rect 4019 3485 4031 3519
rect 3973 3479 4031 3485
rect 4065 3519 4123 3525
rect 4065 3485 4077 3519
rect 4111 3516 4123 3519
rect 4154 3516 4160 3528
rect 4111 3488 4160 3516
rect 4111 3485 4123 3488
rect 4065 3479 4123 3485
rect 2516 3448 2544 3479
rect 4154 3476 4160 3488
rect 4212 3476 4218 3528
rect 4249 3519 4307 3525
rect 4249 3485 4261 3519
rect 4295 3516 4307 3519
rect 4522 3516 4528 3528
rect 4295 3488 4528 3516
rect 4295 3485 4307 3488
rect 4249 3479 4307 3485
rect 4264 3448 4292 3479
rect 4522 3476 4528 3488
rect 4580 3476 4586 3528
rect 5552 3525 5580 3556
rect 5537 3519 5595 3525
rect 5537 3485 5549 3519
rect 5583 3485 5595 3519
rect 5736 3516 5764 3615
rect 5997 3519 6055 3525
rect 5997 3516 6009 3519
rect 5736 3488 6009 3516
rect 5537 3479 5595 3485
rect 5997 3485 6009 3488
rect 6043 3485 6055 3519
rect 5997 3479 6055 3485
rect 2516 3420 4292 3448
rect 4433 3451 4491 3457
rect 4433 3417 4445 3451
rect 4479 3448 4491 3451
rect 4893 3451 4951 3457
rect 4893 3448 4905 3451
rect 4479 3420 4905 3448
rect 4479 3417 4491 3420
rect 4433 3411 4491 3417
rect 4893 3417 4905 3420
rect 4939 3417 4951 3451
rect 4893 3411 4951 3417
rect 3418 3340 3424 3392
rect 3476 3340 3482 3392
rect 6178 3340 6184 3392
rect 6236 3340 6242 3392
rect 1104 3290 6750 3312
rect 1104 3238 2299 3290
rect 2351 3238 2363 3290
rect 2415 3238 2427 3290
rect 2479 3238 2491 3290
rect 2543 3238 2555 3290
rect 2607 3238 3678 3290
rect 3730 3238 3742 3290
rect 3794 3238 3806 3290
rect 3858 3238 3870 3290
rect 3922 3238 3934 3290
rect 3986 3238 5057 3290
rect 5109 3238 5121 3290
rect 5173 3238 5185 3290
rect 5237 3238 5249 3290
rect 5301 3238 5313 3290
rect 5365 3238 6436 3290
rect 6488 3238 6500 3290
rect 6552 3238 6564 3290
rect 6616 3238 6628 3290
rect 6680 3238 6692 3290
rect 6744 3238 6750 3290
rect 1104 3216 6750 3238
rect 3053 3179 3111 3185
rect 3053 3145 3065 3179
rect 3099 3176 3111 3179
rect 3142 3176 3148 3188
rect 3099 3148 3148 3176
rect 3099 3145 3111 3148
rect 3053 3139 3111 3145
rect 3142 3136 3148 3148
rect 3200 3136 3206 3188
rect 4617 3179 4675 3185
rect 4617 3145 4629 3179
rect 4663 3176 4675 3179
rect 4982 3176 4988 3188
rect 4663 3148 4988 3176
rect 4663 3145 4675 3148
rect 4617 3139 4675 3145
rect 4982 3136 4988 3148
rect 5040 3136 5046 3188
rect 2976 3080 4476 3108
rect 2976 3049 3004 3080
rect 2961 3043 3019 3049
rect 2961 3009 2973 3043
rect 3007 3009 3019 3043
rect 2961 3003 3019 3009
rect 3145 3043 3203 3049
rect 3145 3009 3157 3043
rect 3191 3040 3203 3043
rect 4154 3040 4160 3052
rect 3191 3012 4160 3040
rect 3191 3009 3203 3012
rect 3145 3003 3203 3009
rect 4154 3000 4160 3012
rect 4212 3000 4218 3052
rect 4338 3000 4344 3052
rect 4396 3000 4402 3052
rect 4448 3049 4476 3080
rect 4433 3043 4491 3049
rect 4433 3009 4445 3043
rect 4479 3040 4491 3043
rect 4522 3040 4528 3052
rect 4479 3012 4528 3040
rect 4479 3009 4491 3012
rect 4433 3003 4491 3009
rect 4522 3000 4528 3012
rect 4580 3040 4586 3052
rect 4798 3040 4804 3052
rect 4580 3012 4804 3040
rect 4580 3000 4586 3012
rect 4798 3000 4804 3012
rect 4856 3000 4862 3052
rect 3510 2796 3516 2848
rect 3568 2836 3574 2848
rect 4062 2836 4068 2848
rect 3568 2808 4068 2836
rect 3568 2796 3574 2808
rect 4062 2796 4068 2808
rect 4120 2836 4126 2848
rect 4157 2839 4215 2845
rect 4157 2836 4169 2839
rect 4120 2808 4169 2836
rect 4120 2796 4126 2808
rect 4157 2805 4169 2808
rect 4203 2805 4215 2839
rect 4157 2799 4215 2805
rect 1104 2746 6624 2768
rect 1104 2694 1639 2746
rect 1691 2694 1703 2746
rect 1755 2694 1767 2746
rect 1819 2694 1831 2746
rect 1883 2694 1895 2746
rect 1947 2694 3018 2746
rect 3070 2694 3082 2746
rect 3134 2694 3146 2746
rect 3198 2694 3210 2746
rect 3262 2694 3274 2746
rect 3326 2694 4397 2746
rect 4449 2694 4461 2746
rect 4513 2694 4525 2746
rect 4577 2694 4589 2746
rect 4641 2694 4653 2746
rect 4705 2694 5776 2746
rect 5828 2694 5840 2746
rect 5892 2694 5904 2746
rect 5956 2694 5968 2746
rect 6020 2694 6032 2746
rect 6084 2694 6624 2746
rect 1104 2672 6624 2694
rect 3510 2592 3516 2644
rect 3568 2592 3574 2644
rect 4617 2635 4675 2641
rect 4617 2601 4629 2635
rect 4663 2632 4675 2635
rect 4798 2632 4804 2644
rect 4663 2604 4804 2632
rect 4663 2601 4675 2604
rect 4617 2595 4675 2601
rect 4798 2592 4804 2604
rect 4856 2592 4862 2644
rect 2866 2388 2872 2440
rect 2924 2428 2930 2440
rect 2961 2431 3019 2437
rect 2961 2428 2973 2431
rect 2924 2400 2973 2428
rect 2924 2388 2930 2400
rect 2961 2397 2973 2400
rect 3007 2397 3019 2431
rect 2961 2391 3019 2397
rect 3234 2388 3240 2440
rect 3292 2428 3298 2440
rect 3329 2431 3387 2437
rect 3329 2428 3341 2431
rect 3292 2400 3341 2428
rect 3292 2388 3298 2400
rect 3329 2397 3341 2400
rect 3375 2397 3387 2431
rect 3329 2391 3387 2397
rect 3418 2388 3424 2440
rect 3476 2428 3482 2440
rect 3973 2431 4031 2437
rect 3973 2428 3985 2431
rect 3476 2400 3985 2428
rect 3476 2388 3482 2400
rect 3973 2397 3985 2400
rect 4019 2397 4031 2431
rect 3973 2391 4031 2397
rect 4522 2388 4528 2440
rect 4580 2428 4586 2440
rect 4801 2431 4859 2437
rect 4801 2428 4813 2431
rect 4580 2400 4813 2428
rect 4580 2388 4586 2400
rect 4801 2397 4813 2400
rect 4847 2397 4859 2431
rect 4801 2391 4859 2397
rect 2682 2252 2688 2304
rect 2740 2292 2746 2304
rect 2777 2295 2835 2301
rect 2777 2292 2789 2295
rect 2740 2264 2789 2292
rect 2740 2252 2746 2264
rect 2777 2261 2789 2264
rect 2823 2261 2835 2295
rect 2777 2255 2835 2261
rect 4062 2252 4068 2304
rect 4120 2292 4126 2304
rect 4157 2295 4215 2301
rect 4157 2292 4169 2295
rect 4120 2264 4169 2292
rect 4120 2252 4126 2264
rect 4157 2261 4169 2264
rect 4203 2261 4215 2295
rect 4157 2255 4215 2261
rect 1104 2202 6750 2224
rect 1104 2150 2299 2202
rect 2351 2150 2363 2202
rect 2415 2150 2427 2202
rect 2479 2150 2491 2202
rect 2543 2150 2555 2202
rect 2607 2150 3678 2202
rect 3730 2150 3742 2202
rect 3794 2150 3806 2202
rect 3858 2150 3870 2202
rect 3922 2150 3934 2202
rect 3986 2150 5057 2202
rect 5109 2150 5121 2202
rect 5173 2150 5185 2202
rect 5237 2150 5249 2202
rect 5301 2150 5313 2202
rect 5365 2150 6436 2202
rect 6488 2150 6500 2202
rect 6552 2150 6564 2202
rect 6616 2150 6628 2202
rect 6680 2150 6692 2202
rect 6744 2150 6750 2202
rect 1104 2128 6750 2150
<< via1 >>
rect 2299 7590 2351 7642
rect 2363 7590 2415 7642
rect 2427 7590 2479 7642
rect 2491 7590 2543 7642
rect 2555 7590 2607 7642
rect 3678 7590 3730 7642
rect 3742 7590 3794 7642
rect 3806 7590 3858 7642
rect 3870 7590 3922 7642
rect 3934 7590 3986 7642
rect 5057 7590 5109 7642
rect 5121 7590 5173 7642
rect 5185 7590 5237 7642
rect 5249 7590 5301 7642
rect 5313 7590 5365 7642
rect 6436 7590 6488 7642
rect 6500 7590 6552 7642
rect 6564 7590 6616 7642
rect 6628 7590 6680 7642
rect 6692 7590 6744 7642
rect 4068 7488 4120 7540
rect 4804 7531 4856 7540
rect 4804 7497 4813 7531
rect 4813 7497 4847 7531
rect 4847 7497 4856 7531
rect 4804 7488 4856 7497
rect 848 7352 900 7404
rect 1492 7352 1544 7404
rect 2688 7395 2740 7404
rect 2688 7361 2697 7395
rect 2697 7361 2731 7395
rect 2731 7361 2740 7395
rect 2688 7352 2740 7361
rect 3332 7395 3384 7404
rect 3332 7361 3341 7395
rect 3341 7361 3375 7395
rect 3375 7361 3384 7395
rect 3332 7352 3384 7361
rect 4068 7395 4120 7404
rect 4068 7361 4077 7395
rect 4077 7361 4111 7395
rect 4111 7361 4120 7395
rect 4068 7352 4120 7361
rect 4804 7352 4856 7404
rect 1400 7148 1452 7200
rect 2044 7148 2096 7200
rect 2872 7191 2924 7200
rect 2872 7157 2881 7191
rect 2881 7157 2915 7191
rect 2915 7157 2924 7191
rect 2872 7148 2924 7157
rect 3516 7191 3568 7200
rect 3516 7157 3525 7191
rect 3525 7157 3559 7191
rect 3559 7157 3568 7191
rect 3516 7148 3568 7157
rect 1639 7046 1691 7098
rect 1703 7046 1755 7098
rect 1767 7046 1819 7098
rect 1831 7046 1883 7098
rect 1895 7046 1947 7098
rect 3018 7046 3070 7098
rect 3082 7046 3134 7098
rect 3146 7046 3198 7098
rect 3210 7046 3262 7098
rect 3274 7046 3326 7098
rect 4397 7046 4449 7098
rect 4461 7046 4513 7098
rect 4525 7046 4577 7098
rect 4589 7046 4641 7098
rect 4653 7046 4705 7098
rect 5776 7046 5828 7098
rect 5840 7046 5892 7098
rect 5904 7046 5956 7098
rect 5968 7046 6020 7098
rect 6032 7046 6084 7098
rect 4804 6944 4856 6996
rect 4620 6740 4672 6792
rect 2299 6502 2351 6554
rect 2363 6502 2415 6554
rect 2427 6502 2479 6554
rect 2491 6502 2543 6554
rect 2555 6502 2607 6554
rect 3678 6502 3730 6554
rect 3742 6502 3794 6554
rect 3806 6502 3858 6554
rect 3870 6502 3922 6554
rect 3934 6502 3986 6554
rect 5057 6502 5109 6554
rect 5121 6502 5173 6554
rect 5185 6502 5237 6554
rect 5249 6502 5301 6554
rect 5313 6502 5365 6554
rect 6436 6502 6488 6554
rect 6500 6502 6552 6554
rect 6564 6502 6616 6554
rect 6628 6502 6680 6554
rect 6692 6502 6744 6554
rect 1400 6196 1452 6248
rect 2044 6264 2096 6316
rect 2688 6332 2740 6384
rect 2872 6264 2924 6316
rect 3516 6400 3568 6452
rect 4068 6400 4120 6452
rect 4620 6443 4672 6452
rect 4620 6409 4629 6443
rect 4629 6409 4663 6443
rect 4663 6409 4672 6443
rect 4620 6400 4672 6409
rect 4160 6239 4212 6248
rect 4160 6205 4169 6239
rect 4169 6205 4203 6239
rect 4203 6205 4212 6239
rect 4160 6196 4212 6205
rect 2872 6128 2924 6180
rect 1492 6103 1544 6112
rect 1492 6069 1501 6103
rect 1501 6069 1535 6103
rect 1535 6069 1544 6103
rect 1492 6060 1544 6069
rect 2136 6103 2188 6112
rect 2136 6069 2145 6103
rect 2145 6069 2179 6103
rect 2179 6069 2188 6103
rect 2136 6060 2188 6069
rect 2596 6103 2648 6112
rect 2596 6069 2605 6103
rect 2605 6069 2639 6103
rect 2639 6069 2648 6103
rect 2596 6060 2648 6069
rect 3424 6128 3476 6180
rect 4160 6060 4212 6112
rect 1639 5958 1691 6010
rect 1703 5958 1755 6010
rect 1767 5958 1819 6010
rect 1831 5958 1883 6010
rect 1895 5958 1947 6010
rect 3018 5958 3070 6010
rect 3082 5958 3134 6010
rect 3146 5958 3198 6010
rect 3210 5958 3262 6010
rect 3274 5958 3326 6010
rect 4397 5958 4449 6010
rect 4461 5958 4513 6010
rect 4525 5958 4577 6010
rect 4589 5958 4641 6010
rect 4653 5958 4705 6010
rect 5776 5958 5828 6010
rect 5840 5958 5892 6010
rect 5904 5958 5956 6010
rect 5968 5958 6020 6010
rect 6032 5958 6084 6010
rect 1216 5856 1268 5908
rect 3424 5856 3476 5908
rect 2872 5788 2924 5840
rect 1492 5720 1544 5772
rect 2596 5652 2648 5704
rect 2136 5584 2188 5636
rect 2688 5584 2740 5636
rect 6276 5695 6328 5704
rect 6276 5661 6285 5695
rect 6285 5661 6319 5695
rect 6319 5661 6328 5695
rect 6276 5652 6328 5661
rect 1952 5559 2004 5568
rect 1952 5525 1961 5559
rect 1961 5525 1995 5559
rect 1995 5525 2004 5559
rect 1952 5516 2004 5525
rect 5448 5516 5500 5568
rect 2299 5414 2351 5466
rect 2363 5414 2415 5466
rect 2427 5414 2479 5466
rect 2491 5414 2543 5466
rect 2555 5414 2607 5466
rect 3678 5414 3730 5466
rect 3742 5414 3794 5466
rect 3806 5414 3858 5466
rect 3870 5414 3922 5466
rect 3934 5414 3986 5466
rect 5057 5414 5109 5466
rect 5121 5414 5173 5466
rect 5185 5414 5237 5466
rect 5249 5414 5301 5466
rect 5313 5414 5365 5466
rect 6436 5414 6488 5466
rect 6500 5414 6552 5466
rect 6564 5414 6616 5466
rect 6628 5414 6680 5466
rect 6692 5414 6744 5466
rect 5448 5176 5500 5228
rect 4988 5108 5040 5160
rect 6184 4972 6236 5024
rect 1639 4870 1691 4922
rect 1703 4870 1755 4922
rect 1767 4870 1819 4922
rect 1831 4870 1883 4922
rect 1895 4870 1947 4922
rect 3018 4870 3070 4922
rect 3082 4870 3134 4922
rect 3146 4870 3198 4922
rect 3210 4870 3262 4922
rect 3274 4870 3326 4922
rect 4397 4870 4449 4922
rect 4461 4870 4513 4922
rect 4525 4870 4577 4922
rect 4589 4870 4641 4922
rect 4653 4870 4705 4922
rect 5776 4870 5828 4922
rect 5840 4870 5892 4922
rect 5904 4870 5956 4922
rect 5968 4870 6020 4922
rect 6032 4870 6084 4922
rect 6276 4607 6328 4616
rect 6276 4573 6285 4607
rect 6285 4573 6319 4607
rect 6319 4573 6328 4607
rect 6276 4564 6328 4573
rect 4804 4428 4856 4480
rect 2299 4326 2351 4378
rect 2363 4326 2415 4378
rect 2427 4326 2479 4378
rect 2491 4326 2543 4378
rect 2555 4326 2607 4378
rect 3678 4326 3730 4378
rect 3742 4326 3794 4378
rect 3806 4326 3858 4378
rect 3870 4326 3922 4378
rect 3934 4326 3986 4378
rect 5057 4326 5109 4378
rect 5121 4326 5173 4378
rect 5185 4326 5237 4378
rect 5249 4326 5301 4378
rect 5313 4326 5365 4378
rect 6436 4326 6488 4378
rect 6500 4326 6552 4378
rect 6564 4326 6616 4378
rect 6628 4326 6680 4378
rect 6692 4326 6744 4378
rect 2780 4088 2832 4140
rect 3424 4088 3476 4140
rect 2872 3927 2924 3936
rect 2872 3893 2881 3927
rect 2881 3893 2915 3927
rect 2915 3893 2924 3927
rect 2872 3884 2924 3893
rect 1639 3782 1691 3834
rect 1703 3782 1755 3834
rect 1767 3782 1819 3834
rect 1831 3782 1883 3834
rect 1895 3782 1947 3834
rect 3018 3782 3070 3834
rect 3082 3782 3134 3834
rect 3146 3782 3198 3834
rect 3210 3782 3262 3834
rect 3274 3782 3326 3834
rect 4397 3782 4449 3834
rect 4461 3782 4513 3834
rect 4525 3782 4577 3834
rect 4589 3782 4641 3834
rect 4653 3782 4705 3834
rect 5776 3782 5828 3834
rect 5840 3782 5892 3834
rect 5904 3782 5956 3834
rect 5968 3782 6020 3834
rect 6032 3782 6084 3834
rect 2780 3723 2832 3732
rect 2780 3689 2789 3723
rect 2789 3689 2823 3723
rect 2823 3689 2832 3723
rect 2780 3680 2832 3689
rect 4252 3680 4304 3732
rect 4068 3612 4120 3664
rect 4988 3612 5040 3664
rect 3148 3587 3200 3596
rect 3148 3553 3157 3587
rect 3157 3553 3191 3587
rect 3191 3553 3200 3587
rect 3148 3544 3200 3553
rect 3424 3544 3476 3596
rect 4344 3544 4396 3596
rect 4804 3544 4856 3596
rect 4160 3476 4212 3528
rect 4528 3476 4580 3528
rect 3424 3383 3476 3392
rect 3424 3349 3433 3383
rect 3433 3349 3467 3383
rect 3467 3349 3476 3383
rect 3424 3340 3476 3349
rect 6184 3383 6236 3392
rect 6184 3349 6193 3383
rect 6193 3349 6227 3383
rect 6227 3349 6236 3383
rect 6184 3340 6236 3349
rect 2299 3238 2351 3290
rect 2363 3238 2415 3290
rect 2427 3238 2479 3290
rect 2491 3238 2543 3290
rect 2555 3238 2607 3290
rect 3678 3238 3730 3290
rect 3742 3238 3794 3290
rect 3806 3238 3858 3290
rect 3870 3238 3922 3290
rect 3934 3238 3986 3290
rect 5057 3238 5109 3290
rect 5121 3238 5173 3290
rect 5185 3238 5237 3290
rect 5249 3238 5301 3290
rect 5313 3238 5365 3290
rect 6436 3238 6488 3290
rect 6500 3238 6552 3290
rect 6564 3238 6616 3290
rect 6628 3238 6680 3290
rect 6692 3238 6744 3290
rect 3148 3136 3200 3188
rect 4988 3136 5040 3188
rect 4160 3043 4212 3052
rect 4160 3009 4169 3043
rect 4169 3009 4203 3043
rect 4203 3009 4212 3043
rect 4160 3000 4212 3009
rect 4344 3043 4396 3052
rect 4344 3009 4353 3043
rect 4353 3009 4387 3043
rect 4387 3009 4396 3043
rect 4344 3000 4396 3009
rect 4528 3000 4580 3052
rect 4804 3000 4856 3052
rect 3516 2796 3568 2848
rect 4068 2796 4120 2848
rect 1639 2694 1691 2746
rect 1703 2694 1755 2746
rect 1767 2694 1819 2746
rect 1831 2694 1883 2746
rect 1895 2694 1947 2746
rect 3018 2694 3070 2746
rect 3082 2694 3134 2746
rect 3146 2694 3198 2746
rect 3210 2694 3262 2746
rect 3274 2694 3326 2746
rect 4397 2694 4449 2746
rect 4461 2694 4513 2746
rect 4525 2694 4577 2746
rect 4589 2694 4641 2746
rect 4653 2694 4705 2746
rect 5776 2694 5828 2746
rect 5840 2694 5892 2746
rect 5904 2694 5956 2746
rect 5968 2694 6020 2746
rect 6032 2694 6084 2746
rect 3516 2635 3568 2644
rect 3516 2601 3525 2635
rect 3525 2601 3559 2635
rect 3559 2601 3568 2635
rect 3516 2592 3568 2601
rect 4804 2592 4856 2644
rect 2872 2388 2924 2440
rect 3240 2388 3292 2440
rect 3424 2388 3476 2440
rect 4528 2388 4580 2440
rect 2688 2252 2740 2304
rect 4068 2252 4120 2304
rect 2299 2150 2351 2202
rect 2363 2150 2415 2202
rect 2427 2150 2479 2202
rect 2491 2150 2543 2202
rect 2555 2150 2607 2202
rect 3678 2150 3730 2202
rect 3742 2150 3794 2202
rect 3806 2150 3858 2202
rect 3870 2150 3922 2202
rect 3934 2150 3986 2202
rect 5057 2150 5109 2202
rect 5121 2150 5173 2202
rect 5185 2150 5237 2202
rect 5249 2150 5301 2202
rect 5313 2150 5365 2202
rect 6436 2150 6488 2202
rect 6500 2150 6552 2202
rect 6564 2150 6616 2202
rect 6628 2150 6680 2202
rect 6692 2150 6744 2202
<< metal2 >>
rect 2594 9194 2650 9877
rect 3238 9194 3294 9877
rect 3882 9194 3938 9877
rect 4526 9194 4582 9877
rect 2594 9166 2728 9194
rect 2594 9077 2650 9166
rect 2299 7644 2607 7653
rect 2299 7642 2305 7644
rect 2361 7642 2385 7644
rect 2441 7642 2465 7644
rect 2521 7642 2545 7644
rect 2601 7642 2607 7644
rect 2361 7590 2363 7642
rect 2543 7590 2545 7642
rect 2299 7588 2305 7590
rect 2361 7588 2385 7590
rect 2441 7588 2465 7590
rect 2521 7588 2545 7590
rect 2601 7588 2607 7590
rect 2299 7579 2607 7588
rect 846 7440 902 7449
rect 2700 7410 2728 9166
rect 3238 9166 3372 9194
rect 3238 9077 3294 9166
rect 3344 7410 3372 9166
rect 3882 9166 4108 9194
rect 3882 9077 3938 9166
rect 3678 7644 3986 7653
rect 3678 7642 3684 7644
rect 3740 7642 3764 7644
rect 3820 7642 3844 7644
rect 3900 7642 3924 7644
rect 3980 7642 3986 7644
rect 3740 7590 3742 7642
rect 3922 7590 3924 7642
rect 3678 7588 3684 7590
rect 3740 7588 3764 7590
rect 3820 7588 3844 7590
rect 3900 7588 3924 7590
rect 3980 7588 3986 7590
rect 3678 7579 3986 7588
rect 4080 7546 4108 9166
rect 4526 9166 4844 9194
rect 4526 9077 4582 9166
rect 4816 7546 4844 9166
rect 5057 7644 5365 7653
rect 5057 7642 5063 7644
rect 5119 7642 5143 7644
rect 5199 7642 5223 7644
rect 5279 7642 5303 7644
rect 5359 7642 5365 7644
rect 5119 7590 5121 7642
rect 5301 7590 5303 7642
rect 5057 7588 5063 7590
rect 5119 7588 5143 7590
rect 5199 7588 5223 7590
rect 5279 7588 5303 7590
rect 5359 7588 5365 7590
rect 5057 7579 5365 7588
rect 6436 7644 6744 7653
rect 6436 7642 6442 7644
rect 6498 7642 6522 7644
rect 6578 7642 6602 7644
rect 6658 7642 6682 7644
rect 6738 7642 6744 7644
rect 6498 7590 6500 7642
rect 6680 7590 6682 7642
rect 6436 7588 6442 7590
rect 6498 7588 6522 7590
rect 6578 7588 6602 7590
rect 6658 7588 6682 7590
rect 6738 7588 6744 7590
rect 6436 7579 6744 7588
rect 4068 7540 4120 7546
rect 4068 7482 4120 7488
rect 4804 7540 4856 7546
rect 4804 7482 4856 7488
rect 846 7375 848 7384
rect 900 7375 902 7384
rect 1492 7404 1544 7410
rect 848 7346 900 7352
rect 1492 7346 1544 7352
rect 2688 7404 2740 7410
rect 2688 7346 2740 7352
rect 3332 7404 3384 7410
rect 3332 7346 3384 7352
rect 4068 7404 4120 7410
rect 4068 7346 4120 7352
rect 4804 7404 4856 7410
rect 4804 7346 4856 7352
rect 1400 7200 1452 7206
rect 1400 7142 1452 7148
rect 1412 6254 1440 7142
rect 1504 6905 1532 7346
rect 2044 7200 2096 7206
rect 2044 7142 2096 7148
rect 2872 7200 2924 7206
rect 2872 7142 2924 7148
rect 3516 7200 3568 7206
rect 3516 7142 3568 7148
rect 1639 7100 1947 7109
rect 1639 7098 1645 7100
rect 1701 7098 1725 7100
rect 1781 7098 1805 7100
rect 1861 7098 1885 7100
rect 1941 7098 1947 7100
rect 1701 7046 1703 7098
rect 1883 7046 1885 7098
rect 1639 7044 1645 7046
rect 1701 7044 1725 7046
rect 1781 7044 1805 7046
rect 1861 7044 1885 7046
rect 1941 7044 1947 7046
rect 1639 7035 1947 7044
rect 1490 6896 1546 6905
rect 1490 6831 1546 6840
rect 2056 6322 2084 7142
rect 2299 6556 2607 6565
rect 2299 6554 2305 6556
rect 2361 6554 2385 6556
rect 2441 6554 2465 6556
rect 2521 6554 2545 6556
rect 2601 6554 2607 6556
rect 2361 6502 2363 6554
rect 2543 6502 2545 6554
rect 2299 6500 2305 6502
rect 2361 6500 2385 6502
rect 2441 6500 2465 6502
rect 2521 6500 2545 6502
rect 2601 6500 2607 6502
rect 2299 6491 2607 6500
rect 2688 6384 2740 6390
rect 2688 6326 2740 6332
rect 2044 6316 2096 6322
rect 2044 6258 2096 6264
rect 1400 6248 1452 6254
rect 1214 6216 1270 6225
rect 1400 6190 1452 6196
rect 1214 6151 1270 6160
rect 1228 5914 1256 6151
rect 1492 6112 1544 6118
rect 1492 6054 1544 6060
rect 2136 6112 2188 6118
rect 2136 6054 2188 6060
rect 2596 6112 2648 6118
rect 2596 6054 2648 6060
rect 1216 5908 1268 5914
rect 1216 5850 1268 5856
rect 1504 5778 1532 6054
rect 1639 6012 1947 6021
rect 1639 6010 1645 6012
rect 1701 6010 1725 6012
rect 1781 6010 1805 6012
rect 1861 6010 1885 6012
rect 1941 6010 1947 6012
rect 1701 5958 1703 6010
rect 1883 5958 1885 6010
rect 1639 5956 1645 5958
rect 1701 5956 1725 5958
rect 1781 5956 1805 5958
rect 1861 5956 1885 5958
rect 1941 5956 1947 5958
rect 1639 5947 1947 5956
rect 1492 5772 1544 5778
rect 1492 5714 1544 5720
rect 2148 5642 2176 6054
rect 2608 5710 2636 6054
rect 2596 5704 2648 5710
rect 2596 5646 2648 5652
rect 2700 5642 2728 6326
rect 2884 6322 2912 7142
rect 3018 7100 3326 7109
rect 3018 7098 3024 7100
rect 3080 7098 3104 7100
rect 3160 7098 3184 7100
rect 3240 7098 3264 7100
rect 3320 7098 3326 7100
rect 3080 7046 3082 7098
rect 3262 7046 3264 7098
rect 3018 7044 3024 7046
rect 3080 7044 3104 7046
rect 3160 7044 3184 7046
rect 3240 7044 3264 7046
rect 3320 7044 3326 7046
rect 3018 7035 3326 7044
rect 3528 6458 3556 7142
rect 3678 6556 3986 6565
rect 3678 6554 3684 6556
rect 3740 6554 3764 6556
rect 3820 6554 3844 6556
rect 3900 6554 3924 6556
rect 3980 6554 3986 6556
rect 3740 6502 3742 6554
rect 3922 6502 3924 6554
rect 3678 6500 3684 6502
rect 3740 6500 3764 6502
rect 3820 6500 3844 6502
rect 3900 6500 3924 6502
rect 3980 6500 3986 6502
rect 3678 6491 3986 6500
rect 4080 6458 4108 7346
rect 4397 7100 4705 7109
rect 4397 7098 4403 7100
rect 4459 7098 4483 7100
rect 4539 7098 4563 7100
rect 4619 7098 4643 7100
rect 4699 7098 4705 7100
rect 4459 7046 4461 7098
rect 4641 7046 4643 7098
rect 4397 7044 4403 7046
rect 4459 7044 4483 7046
rect 4539 7044 4563 7046
rect 4619 7044 4643 7046
rect 4699 7044 4705 7046
rect 4397 7035 4705 7044
rect 4816 7002 4844 7346
rect 5776 7100 6084 7109
rect 5776 7098 5782 7100
rect 5838 7098 5862 7100
rect 5918 7098 5942 7100
rect 5998 7098 6022 7100
rect 6078 7098 6084 7100
rect 5838 7046 5840 7098
rect 6020 7046 6022 7098
rect 5776 7044 5782 7046
rect 5838 7044 5862 7046
rect 5918 7044 5942 7046
rect 5998 7044 6022 7046
rect 6078 7044 6084 7046
rect 5776 7035 6084 7044
rect 4804 6996 4856 7002
rect 4804 6938 4856 6944
rect 4620 6792 4672 6798
rect 4620 6734 4672 6740
rect 4632 6458 4660 6734
rect 5057 6556 5365 6565
rect 5057 6554 5063 6556
rect 5119 6554 5143 6556
rect 5199 6554 5223 6556
rect 5279 6554 5303 6556
rect 5359 6554 5365 6556
rect 5119 6502 5121 6554
rect 5301 6502 5303 6554
rect 5057 6500 5063 6502
rect 5119 6500 5143 6502
rect 5199 6500 5223 6502
rect 5279 6500 5303 6502
rect 5359 6500 5365 6502
rect 5057 6491 5365 6500
rect 6436 6556 6744 6565
rect 6436 6554 6442 6556
rect 6498 6554 6522 6556
rect 6578 6554 6602 6556
rect 6658 6554 6682 6556
rect 6738 6554 6744 6556
rect 6498 6502 6500 6554
rect 6680 6502 6682 6554
rect 6436 6500 6442 6502
rect 6498 6500 6522 6502
rect 6578 6500 6602 6502
rect 6658 6500 6682 6502
rect 6738 6500 6744 6502
rect 6436 6491 6744 6500
rect 3516 6452 3568 6458
rect 3516 6394 3568 6400
rect 4068 6452 4120 6458
rect 4068 6394 4120 6400
rect 4620 6452 4672 6458
rect 4620 6394 4672 6400
rect 2872 6316 2924 6322
rect 2872 6258 2924 6264
rect 2884 6186 2912 6258
rect 4160 6248 4212 6254
rect 4160 6190 4212 6196
rect 2872 6180 2924 6186
rect 2872 6122 2924 6128
rect 3424 6180 3476 6186
rect 3424 6122 3476 6128
rect 2884 5846 2912 6122
rect 3018 6012 3326 6021
rect 3018 6010 3024 6012
rect 3080 6010 3104 6012
rect 3160 6010 3184 6012
rect 3240 6010 3264 6012
rect 3320 6010 3326 6012
rect 3080 5958 3082 6010
rect 3262 5958 3264 6010
rect 3018 5956 3024 5958
rect 3080 5956 3104 5958
rect 3160 5956 3184 5958
rect 3240 5956 3264 5958
rect 3320 5956 3326 5958
rect 3018 5947 3326 5956
rect 3436 5914 3464 6122
rect 4172 6118 4200 6190
rect 4160 6112 4212 6118
rect 4160 6054 4212 6060
rect 3424 5908 3476 5914
rect 3424 5850 3476 5856
rect 2872 5840 2924 5846
rect 2872 5782 2924 5788
rect 2136 5636 2188 5642
rect 2136 5578 2188 5584
rect 2688 5636 2740 5642
rect 2688 5578 2740 5584
rect 1952 5568 2004 5574
rect 1950 5536 1952 5545
rect 2004 5536 2006 5545
rect 1950 5471 2006 5480
rect 2299 5468 2607 5477
rect 2299 5466 2305 5468
rect 2361 5466 2385 5468
rect 2441 5466 2465 5468
rect 2521 5466 2545 5468
rect 2601 5466 2607 5468
rect 2361 5414 2363 5466
rect 2543 5414 2545 5466
rect 2299 5412 2305 5414
rect 2361 5412 2385 5414
rect 2441 5412 2465 5414
rect 2521 5412 2545 5414
rect 2601 5412 2607 5414
rect 2299 5403 2607 5412
rect 3678 5468 3986 5477
rect 3678 5466 3684 5468
rect 3740 5466 3764 5468
rect 3820 5466 3844 5468
rect 3900 5466 3924 5468
rect 3980 5466 3986 5468
rect 3740 5414 3742 5466
rect 3922 5414 3924 5466
rect 3678 5412 3684 5414
rect 3740 5412 3764 5414
rect 3820 5412 3844 5414
rect 3900 5412 3924 5414
rect 3980 5412 3986 5414
rect 3678 5403 3986 5412
rect 1639 4924 1947 4933
rect 1639 4922 1645 4924
rect 1701 4922 1725 4924
rect 1781 4922 1805 4924
rect 1861 4922 1885 4924
rect 1941 4922 1947 4924
rect 1701 4870 1703 4922
rect 1883 4870 1885 4922
rect 1639 4868 1645 4870
rect 1701 4868 1725 4870
rect 1781 4868 1805 4870
rect 1861 4868 1885 4870
rect 1941 4868 1947 4870
rect 1639 4859 1947 4868
rect 3018 4924 3326 4933
rect 3018 4922 3024 4924
rect 3080 4922 3104 4924
rect 3160 4922 3184 4924
rect 3240 4922 3264 4924
rect 3320 4922 3326 4924
rect 3080 4870 3082 4922
rect 3262 4870 3264 4922
rect 3018 4868 3024 4870
rect 3080 4868 3104 4870
rect 3160 4868 3184 4870
rect 3240 4868 3264 4870
rect 3320 4868 3326 4870
rect 3018 4859 3326 4868
rect 2299 4380 2607 4389
rect 2299 4378 2305 4380
rect 2361 4378 2385 4380
rect 2441 4378 2465 4380
rect 2521 4378 2545 4380
rect 2601 4378 2607 4380
rect 2361 4326 2363 4378
rect 2543 4326 2545 4378
rect 2299 4324 2305 4326
rect 2361 4324 2385 4326
rect 2441 4324 2465 4326
rect 2521 4324 2545 4326
rect 2601 4324 2607 4326
rect 2299 4315 2607 4324
rect 3678 4380 3986 4389
rect 3678 4378 3684 4380
rect 3740 4378 3764 4380
rect 3820 4378 3844 4380
rect 3900 4378 3924 4380
rect 3980 4378 3986 4380
rect 3740 4326 3742 4378
rect 3922 4326 3924 4378
rect 3678 4324 3684 4326
rect 3740 4324 3764 4326
rect 3820 4324 3844 4326
rect 3900 4324 3924 4326
rect 3980 4324 3986 4326
rect 3678 4315 3986 4324
rect 2780 4140 2832 4146
rect 2780 4082 2832 4088
rect 3424 4140 3476 4146
rect 3424 4082 3476 4088
rect 1639 3836 1947 3845
rect 1639 3834 1645 3836
rect 1701 3834 1725 3836
rect 1781 3834 1805 3836
rect 1861 3834 1885 3836
rect 1941 3834 1947 3836
rect 1701 3782 1703 3834
rect 1883 3782 1885 3834
rect 1639 3780 1645 3782
rect 1701 3780 1725 3782
rect 1781 3780 1805 3782
rect 1861 3780 1885 3782
rect 1941 3780 1947 3782
rect 1639 3771 1947 3780
rect 2792 3738 2820 4082
rect 2872 3936 2924 3942
rect 2872 3878 2924 3884
rect 2780 3732 2832 3738
rect 2780 3674 2832 3680
rect 2299 3292 2607 3301
rect 2299 3290 2305 3292
rect 2361 3290 2385 3292
rect 2441 3290 2465 3292
rect 2521 3290 2545 3292
rect 2601 3290 2607 3292
rect 2361 3238 2363 3290
rect 2543 3238 2545 3290
rect 2299 3236 2305 3238
rect 2361 3236 2385 3238
rect 2441 3236 2465 3238
rect 2521 3236 2545 3238
rect 2601 3236 2607 3238
rect 2299 3227 2607 3236
rect 1639 2748 1947 2757
rect 1639 2746 1645 2748
rect 1701 2746 1725 2748
rect 1781 2746 1805 2748
rect 1861 2746 1885 2748
rect 1941 2746 1947 2748
rect 1701 2694 1703 2746
rect 1883 2694 1885 2746
rect 1639 2692 1645 2694
rect 1701 2692 1725 2694
rect 1781 2692 1805 2694
rect 1861 2692 1885 2694
rect 1941 2692 1947 2694
rect 1639 2683 1947 2692
rect 2884 2446 2912 3878
rect 3018 3836 3326 3845
rect 3018 3834 3024 3836
rect 3080 3834 3104 3836
rect 3160 3834 3184 3836
rect 3240 3834 3264 3836
rect 3320 3834 3326 3836
rect 3080 3782 3082 3834
rect 3262 3782 3264 3834
rect 3018 3780 3024 3782
rect 3080 3780 3104 3782
rect 3160 3780 3184 3782
rect 3240 3780 3264 3782
rect 3320 3780 3326 3782
rect 3018 3771 3326 3780
rect 3436 3602 3464 4082
rect 4172 3754 4200 6054
rect 4397 6012 4705 6021
rect 4397 6010 4403 6012
rect 4459 6010 4483 6012
rect 4539 6010 4563 6012
rect 4619 6010 4643 6012
rect 4699 6010 4705 6012
rect 4459 5958 4461 6010
rect 4641 5958 4643 6010
rect 4397 5956 4403 5958
rect 4459 5956 4483 5958
rect 4539 5956 4563 5958
rect 4619 5956 4643 5958
rect 4699 5956 4705 5958
rect 4397 5947 4705 5956
rect 5776 6012 6084 6021
rect 5776 6010 5782 6012
rect 5838 6010 5862 6012
rect 5918 6010 5942 6012
rect 5998 6010 6022 6012
rect 6078 6010 6084 6012
rect 5838 5958 5840 6010
rect 6020 5958 6022 6010
rect 5776 5956 5782 5958
rect 5838 5956 5862 5958
rect 5918 5956 5942 5958
rect 5998 5956 6022 5958
rect 6078 5956 6084 5958
rect 5776 5947 6084 5956
rect 6274 5808 6330 5817
rect 6274 5743 6330 5752
rect 6288 5710 6316 5743
rect 6276 5704 6328 5710
rect 6276 5646 6328 5652
rect 5448 5568 5500 5574
rect 5448 5510 5500 5516
rect 5057 5468 5365 5477
rect 5057 5466 5063 5468
rect 5119 5466 5143 5468
rect 5199 5466 5223 5468
rect 5279 5466 5303 5468
rect 5359 5466 5365 5468
rect 5119 5414 5121 5466
rect 5301 5414 5303 5466
rect 5057 5412 5063 5414
rect 5119 5412 5143 5414
rect 5199 5412 5223 5414
rect 5279 5412 5303 5414
rect 5359 5412 5365 5414
rect 5057 5403 5365 5412
rect 5460 5234 5488 5510
rect 6436 5468 6744 5477
rect 6436 5466 6442 5468
rect 6498 5466 6522 5468
rect 6578 5466 6602 5468
rect 6658 5466 6682 5468
rect 6738 5466 6744 5468
rect 6498 5414 6500 5466
rect 6680 5414 6682 5466
rect 6436 5412 6442 5414
rect 6498 5412 6522 5414
rect 6578 5412 6602 5414
rect 6658 5412 6682 5414
rect 6738 5412 6744 5414
rect 6436 5403 6744 5412
rect 5448 5228 5500 5234
rect 5448 5170 5500 5176
rect 4988 5160 5040 5166
rect 4988 5102 5040 5108
rect 4397 4924 4705 4933
rect 4397 4922 4403 4924
rect 4459 4922 4483 4924
rect 4539 4922 4563 4924
rect 4619 4922 4643 4924
rect 4699 4922 4705 4924
rect 4459 4870 4461 4922
rect 4641 4870 4643 4922
rect 4397 4868 4403 4870
rect 4459 4868 4483 4870
rect 4539 4868 4563 4870
rect 4619 4868 4643 4870
rect 4699 4868 4705 4870
rect 4397 4859 4705 4868
rect 4804 4480 4856 4486
rect 4804 4422 4856 4428
rect 4397 3836 4705 3845
rect 4397 3834 4403 3836
rect 4459 3834 4483 3836
rect 4539 3834 4563 3836
rect 4619 3834 4643 3836
rect 4699 3834 4705 3836
rect 4459 3782 4461 3834
rect 4641 3782 4643 3834
rect 4397 3780 4403 3782
rect 4459 3780 4483 3782
rect 4539 3780 4563 3782
rect 4619 3780 4643 3782
rect 4699 3780 4705 3782
rect 4397 3771 4705 3780
rect 4172 3738 4292 3754
rect 4172 3732 4304 3738
rect 4172 3726 4252 3732
rect 4068 3664 4120 3670
rect 4068 3606 4120 3612
rect 3148 3596 3200 3602
rect 3148 3538 3200 3544
rect 3424 3596 3476 3602
rect 3424 3538 3476 3544
rect 3160 3194 3188 3538
rect 3424 3392 3476 3398
rect 3424 3334 3476 3340
rect 3148 3188 3200 3194
rect 3148 3130 3200 3136
rect 3018 2748 3326 2757
rect 3018 2746 3024 2748
rect 3080 2746 3104 2748
rect 3160 2746 3184 2748
rect 3240 2746 3264 2748
rect 3320 2746 3326 2748
rect 3080 2694 3082 2746
rect 3262 2694 3264 2746
rect 3018 2692 3024 2694
rect 3080 2692 3104 2694
rect 3160 2692 3184 2694
rect 3240 2692 3264 2694
rect 3320 2692 3326 2694
rect 3018 2683 3326 2692
rect 3436 2446 3464 3334
rect 3678 3292 3986 3301
rect 3678 3290 3684 3292
rect 3740 3290 3764 3292
rect 3820 3290 3844 3292
rect 3900 3290 3924 3292
rect 3980 3290 3986 3292
rect 3740 3238 3742 3290
rect 3922 3238 3924 3290
rect 3678 3236 3684 3238
rect 3740 3236 3764 3238
rect 3820 3236 3844 3238
rect 3900 3236 3924 3238
rect 3980 3236 3986 3238
rect 3678 3227 3986 3236
rect 4080 2854 4108 3606
rect 4172 3534 4200 3726
rect 4252 3674 4304 3680
rect 4816 3602 4844 4422
rect 5000 3670 5028 5102
rect 6184 5024 6236 5030
rect 6184 4966 6236 4972
rect 5776 4924 6084 4933
rect 5776 4922 5782 4924
rect 5838 4922 5862 4924
rect 5918 4922 5942 4924
rect 5998 4922 6022 4924
rect 6078 4922 6084 4924
rect 5838 4870 5840 4922
rect 6020 4870 6022 4922
rect 5776 4868 5782 4870
rect 5838 4868 5862 4870
rect 5918 4868 5942 4870
rect 5998 4868 6022 4870
rect 6078 4868 6084 4870
rect 5776 4859 6084 4868
rect 6196 4865 6224 4966
rect 6182 4856 6238 4865
rect 6182 4791 6238 4800
rect 6276 4616 6328 4622
rect 6276 4558 6328 4564
rect 5057 4380 5365 4389
rect 5057 4378 5063 4380
rect 5119 4378 5143 4380
rect 5199 4378 5223 4380
rect 5279 4378 5303 4380
rect 5359 4378 5365 4380
rect 5119 4326 5121 4378
rect 5301 4326 5303 4378
rect 5057 4324 5063 4326
rect 5119 4324 5143 4326
rect 5199 4324 5223 4326
rect 5279 4324 5303 4326
rect 5359 4324 5365 4326
rect 5057 4315 5365 4324
rect 6288 4185 6316 4558
rect 6436 4380 6744 4389
rect 6436 4378 6442 4380
rect 6498 4378 6522 4380
rect 6578 4378 6602 4380
rect 6658 4378 6682 4380
rect 6738 4378 6744 4380
rect 6498 4326 6500 4378
rect 6680 4326 6682 4378
rect 6436 4324 6442 4326
rect 6498 4324 6522 4326
rect 6578 4324 6602 4326
rect 6658 4324 6682 4326
rect 6738 4324 6744 4326
rect 6436 4315 6744 4324
rect 6274 4176 6330 4185
rect 6274 4111 6330 4120
rect 5776 3836 6084 3845
rect 5776 3834 5782 3836
rect 5838 3834 5862 3836
rect 5918 3834 5942 3836
rect 5998 3834 6022 3836
rect 6078 3834 6084 3836
rect 5838 3782 5840 3834
rect 6020 3782 6022 3834
rect 5776 3780 5782 3782
rect 5838 3780 5862 3782
rect 5918 3780 5942 3782
rect 5998 3780 6022 3782
rect 6078 3780 6084 3782
rect 5776 3771 6084 3780
rect 4988 3664 5040 3670
rect 4988 3606 5040 3612
rect 4344 3596 4396 3602
rect 4344 3538 4396 3544
rect 4804 3596 4856 3602
rect 4804 3538 4856 3544
rect 4160 3528 4212 3534
rect 4160 3470 4212 3476
rect 4172 3058 4200 3470
rect 4356 3058 4384 3538
rect 4528 3528 4580 3534
rect 4528 3470 4580 3476
rect 4540 3058 4568 3470
rect 5000 3194 5028 3606
rect 6182 3496 6238 3505
rect 6182 3431 6238 3440
rect 6196 3398 6224 3431
rect 6184 3392 6236 3398
rect 6184 3334 6236 3340
rect 5057 3292 5365 3301
rect 5057 3290 5063 3292
rect 5119 3290 5143 3292
rect 5199 3290 5223 3292
rect 5279 3290 5303 3292
rect 5359 3290 5365 3292
rect 5119 3238 5121 3290
rect 5301 3238 5303 3290
rect 5057 3236 5063 3238
rect 5119 3236 5143 3238
rect 5199 3236 5223 3238
rect 5279 3236 5303 3238
rect 5359 3236 5365 3238
rect 5057 3227 5365 3236
rect 6436 3292 6744 3301
rect 6436 3290 6442 3292
rect 6498 3290 6522 3292
rect 6578 3290 6602 3292
rect 6658 3290 6682 3292
rect 6738 3290 6744 3292
rect 6498 3238 6500 3290
rect 6680 3238 6682 3290
rect 6436 3236 6442 3238
rect 6498 3236 6522 3238
rect 6578 3236 6602 3238
rect 6658 3236 6682 3238
rect 6738 3236 6744 3238
rect 6436 3227 6744 3236
rect 4988 3188 5040 3194
rect 4988 3130 5040 3136
rect 4160 3052 4212 3058
rect 4160 2994 4212 3000
rect 4344 3052 4396 3058
rect 4344 2994 4396 3000
rect 4528 3052 4580 3058
rect 4528 2994 4580 3000
rect 4804 3052 4856 3058
rect 4804 2994 4856 3000
rect 3516 2848 3568 2854
rect 3516 2790 3568 2796
rect 4068 2848 4120 2854
rect 4068 2790 4120 2796
rect 3528 2650 3556 2790
rect 4397 2748 4705 2757
rect 4397 2746 4403 2748
rect 4459 2746 4483 2748
rect 4539 2746 4563 2748
rect 4619 2746 4643 2748
rect 4699 2746 4705 2748
rect 4459 2694 4461 2746
rect 4641 2694 4643 2746
rect 4397 2692 4403 2694
rect 4459 2692 4483 2694
rect 4539 2692 4563 2694
rect 4619 2692 4643 2694
rect 4699 2692 4705 2694
rect 4397 2683 4705 2692
rect 4816 2650 4844 2994
rect 5776 2748 6084 2757
rect 5776 2746 5782 2748
rect 5838 2746 5862 2748
rect 5918 2746 5942 2748
rect 5998 2746 6022 2748
rect 6078 2746 6084 2748
rect 5838 2694 5840 2746
rect 6020 2694 6022 2746
rect 5776 2692 5782 2694
rect 5838 2692 5862 2694
rect 5918 2692 5942 2694
rect 5998 2692 6022 2694
rect 6078 2692 6084 2694
rect 5776 2683 6084 2692
rect 3516 2644 3568 2650
rect 3516 2586 3568 2592
rect 4804 2644 4856 2650
rect 4804 2586 4856 2592
rect 2872 2440 2924 2446
rect 2872 2382 2924 2388
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 3424 2440 3476 2446
rect 3424 2382 3476 2388
rect 4528 2440 4580 2446
rect 4528 2382 4580 2388
rect 2688 2304 2740 2310
rect 2688 2246 2740 2252
rect 2299 2204 2607 2213
rect 2299 2202 2305 2204
rect 2361 2202 2385 2204
rect 2441 2202 2465 2204
rect 2521 2202 2545 2204
rect 2601 2202 2607 2204
rect 2361 2150 2363 2202
rect 2543 2150 2545 2202
rect 2299 2148 2305 2150
rect 2361 2148 2385 2150
rect 2441 2148 2465 2150
rect 2521 2148 2545 2150
rect 2601 2148 2607 2150
rect 2299 2139 2607 2148
rect 2700 1170 2728 2246
rect 2608 1142 2728 1170
rect 2608 800 2636 1142
rect 3252 800 3280 2382
rect 4068 2304 4120 2310
rect 4068 2246 4120 2252
rect 3678 2204 3986 2213
rect 3678 2202 3684 2204
rect 3740 2202 3764 2204
rect 3820 2202 3844 2204
rect 3900 2202 3924 2204
rect 3980 2202 3986 2204
rect 3740 2150 3742 2202
rect 3922 2150 3924 2202
rect 3678 2148 3684 2150
rect 3740 2148 3764 2150
rect 3820 2148 3844 2150
rect 3900 2148 3924 2150
rect 3980 2148 3986 2150
rect 3678 2139 3986 2148
rect 4080 1170 4108 2246
rect 3896 1142 4108 1170
rect 3896 800 3924 1142
rect 4540 800 4568 2382
rect 5057 2204 5365 2213
rect 5057 2202 5063 2204
rect 5119 2202 5143 2204
rect 5199 2202 5223 2204
rect 5279 2202 5303 2204
rect 5359 2202 5365 2204
rect 5119 2150 5121 2202
rect 5301 2150 5303 2202
rect 5057 2148 5063 2150
rect 5119 2148 5143 2150
rect 5199 2148 5223 2150
rect 5279 2148 5303 2150
rect 5359 2148 5365 2150
rect 5057 2139 5365 2148
rect 6436 2204 6744 2213
rect 6436 2202 6442 2204
rect 6498 2202 6522 2204
rect 6578 2202 6602 2204
rect 6658 2202 6682 2204
rect 6738 2202 6744 2204
rect 6498 2150 6500 2202
rect 6680 2150 6682 2202
rect 6436 2148 6442 2150
rect 6498 2148 6522 2150
rect 6578 2148 6602 2150
rect 6658 2148 6682 2150
rect 6738 2148 6744 2150
rect 6436 2139 6744 2148
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
<< via2 >>
rect 2305 7642 2361 7644
rect 2385 7642 2441 7644
rect 2465 7642 2521 7644
rect 2545 7642 2601 7644
rect 2305 7590 2351 7642
rect 2351 7590 2361 7642
rect 2385 7590 2415 7642
rect 2415 7590 2427 7642
rect 2427 7590 2441 7642
rect 2465 7590 2479 7642
rect 2479 7590 2491 7642
rect 2491 7590 2521 7642
rect 2545 7590 2555 7642
rect 2555 7590 2601 7642
rect 2305 7588 2361 7590
rect 2385 7588 2441 7590
rect 2465 7588 2521 7590
rect 2545 7588 2601 7590
rect 846 7404 902 7440
rect 3684 7642 3740 7644
rect 3764 7642 3820 7644
rect 3844 7642 3900 7644
rect 3924 7642 3980 7644
rect 3684 7590 3730 7642
rect 3730 7590 3740 7642
rect 3764 7590 3794 7642
rect 3794 7590 3806 7642
rect 3806 7590 3820 7642
rect 3844 7590 3858 7642
rect 3858 7590 3870 7642
rect 3870 7590 3900 7642
rect 3924 7590 3934 7642
rect 3934 7590 3980 7642
rect 3684 7588 3740 7590
rect 3764 7588 3820 7590
rect 3844 7588 3900 7590
rect 3924 7588 3980 7590
rect 5063 7642 5119 7644
rect 5143 7642 5199 7644
rect 5223 7642 5279 7644
rect 5303 7642 5359 7644
rect 5063 7590 5109 7642
rect 5109 7590 5119 7642
rect 5143 7590 5173 7642
rect 5173 7590 5185 7642
rect 5185 7590 5199 7642
rect 5223 7590 5237 7642
rect 5237 7590 5249 7642
rect 5249 7590 5279 7642
rect 5303 7590 5313 7642
rect 5313 7590 5359 7642
rect 5063 7588 5119 7590
rect 5143 7588 5199 7590
rect 5223 7588 5279 7590
rect 5303 7588 5359 7590
rect 6442 7642 6498 7644
rect 6522 7642 6578 7644
rect 6602 7642 6658 7644
rect 6682 7642 6738 7644
rect 6442 7590 6488 7642
rect 6488 7590 6498 7642
rect 6522 7590 6552 7642
rect 6552 7590 6564 7642
rect 6564 7590 6578 7642
rect 6602 7590 6616 7642
rect 6616 7590 6628 7642
rect 6628 7590 6658 7642
rect 6682 7590 6692 7642
rect 6692 7590 6738 7642
rect 6442 7588 6498 7590
rect 6522 7588 6578 7590
rect 6602 7588 6658 7590
rect 6682 7588 6738 7590
rect 846 7384 848 7404
rect 848 7384 900 7404
rect 900 7384 902 7404
rect 1645 7098 1701 7100
rect 1725 7098 1781 7100
rect 1805 7098 1861 7100
rect 1885 7098 1941 7100
rect 1645 7046 1691 7098
rect 1691 7046 1701 7098
rect 1725 7046 1755 7098
rect 1755 7046 1767 7098
rect 1767 7046 1781 7098
rect 1805 7046 1819 7098
rect 1819 7046 1831 7098
rect 1831 7046 1861 7098
rect 1885 7046 1895 7098
rect 1895 7046 1941 7098
rect 1645 7044 1701 7046
rect 1725 7044 1781 7046
rect 1805 7044 1861 7046
rect 1885 7044 1941 7046
rect 1490 6840 1546 6896
rect 2305 6554 2361 6556
rect 2385 6554 2441 6556
rect 2465 6554 2521 6556
rect 2545 6554 2601 6556
rect 2305 6502 2351 6554
rect 2351 6502 2361 6554
rect 2385 6502 2415 6554
rect 2415 6502 2427 6554
rect 2427 6502 2441 6554
rect 2465 6502 2479 6554
rect 2479 6502 2491 6554
rect 2491 6502 2521 6554
rect 2545 6502 2555 6554
rect 2555 6502 2601 6554
rect 2305 6500 2361 6502
rect 2385 6500 2441 6502
rect 2465 6500 2521 6502
rect 2545 6500 2601 6502
rect 1214 6160 1270 6216
rect 1645 6010 1701 6012
rect 1725 6010 1781 6012
rect 1805 6010 1861 6012
rect 1885 6010 1941 6012
rect 1645 5958 1691 6010
rect 1691 5958 1701 6010
rect 1725 5958 1755 6010
rect 1755 5958 1767 6010
rect 1767 5958 1781 6010
rect 1805 5958 1819 6010
rect 1819 5958 1831 6010
rect 1831 5958 1861 6010
rect 1885 5958 1895 6010
rect 1895 5958 1941 6010
rect 1645 5956 1701 5958
rect 1725 5956 1781 5958
rect 1805 5956 1861 5958
rect 1885 5956 1941 5958
rect 3024 7098 3080 7100
rect 3104 7098 3160 7100
rect 3184 7098 3240 7100
rect 3264 7098 3320 7100
rect 3024 7046 3070 7098
rect 3070 7046 3080 7098
rect 3104 7046 3134 7098
rect 3134 7046 3146 7098
rect 3146 7046 3160 7098
rect 3184 7046 3198 7098
rect 3198 7046 3210 7098
rect 3210 7046 3240 7098
rect 3264 7046 3274 7098
rect 3274 7046 3320 7098
rect 3024 7044 3080 7046
rect 3104 7044 3160 7046
rect 3184 7044 3240 7046
rect 3264 7044 3320 7046
rect 3684 6554 3740 6556
rect 3764 6554 3820 6556
rect 3844 6554 3900 6556
rect 3924 6554 3980 6556
rect 3684 6502 3730 6554
rect 3730 6502 3740 6554
rect 3764 6502 3794 6554
rect 3794 6502 3806 6554
rect 3806 6502 3820 6554
rect 3844 6502 3858 6554
rect 3858 6502 3870 6554
rect 3870 6502 3900 6554
rect 3924 6502 3934 6554
rect 3934 6502 3980 6554
rect 3684 6500 3740 6502
rect 3764 6500 3820 6502
rect 3844 6500 3900 6502
rect 3924 6500 3980 6502
rect 4403 7098 4459 7100
rect 4483 7098 4539 7100
rect 4563 7098 4619 7100
rect 4643 7098 4699 7100
rect 4403 7046 4449 7098
rect 4449 7046 4459 7098
rect 4483 7046 4513 7098
rect 4513 7046 4525 7098
rect 4525 7046 4539 7098
rect 4563 7046 4577 7098
rect 4577 7046 4589 7098
rect 4589 7046 4619 7098
rect 4643 7046 4653 7098
rect 4653 7046 4699 7098
rect 4403 7044 4459 7046
rect 4483 7044 4539 7046
rect 4563 7044 4619 7046
rect 4643 7044 4699 7046
rect 5782 7098 5838 7100
rect 5862 7098 5918 7100
rect 5942 7098 5998 7100
rect 6022 7098 6078 7100
rect 5782 7046 5828 7098
rect 5828 7046 5838 7098
rect 5862 7046 5892 7098
rect 5892 7046 5904 7098
rect 5904 7046 5918 7098
rect 5942 7046 5956 7098
rect 5956 7046 5968 7098
rect 5968 7046 5998 7098
rect 6022 7046 6032 7098
rect 6032 7046 6078 7098
rect 5782 7044 5838 7046
rect 5862 7044 5918 7046
rect 5942 7044 5998 7046
rect 6022 7044 6078 7046
rect 5063 6554 5119 6556
rect 5143 6554 5199 6556
rect 5223 6554 5279 6556
rect 5303 6554 5359 6556
rect 5063 6502 5109 6554
rect 5109 6502 5119 6554
rect 5143 6502 5173 6554
rect 5173 6502 5185 6554
rect 5185 6502 5199 6554
rect 5223 6502 5237 6554
rect 5237 6502 5249 6554
rect 5249 6502 5279 6554
rect 5303 6502 5313 6554
rect 5313 6502 5359 6554
rect 5063 6500 5119 6502
rect 5143 6500 5199 6502
rect 5223 6500 5279 6502
rect 5303 6500 5359 6502
rect 6442 6554 6498 6556
rect 6522 6554 6578 6556
rect 6602 6554 6658 6556
rect 6682 6554 6738 6556
rect 6442 6502 6488 6554
rect 6488 6502 6498 6554
rect 6522 6502 6552 6554
rect 6552 6502 6564 6554
rect 6564 6502 6578 6554
rect 6602 6502 6616 6554
rect 6616 6502 6628 6554
rect 6628 6502 6658 6554
rect 6682 6502 6692 6554
rect 6692 6502 6738 6554
rect 6442 6500 6498 6502
rect 6522 6500 6578 6502
rect 6602 6500 6658 6502
rect 6682 6500 6738 6502
rect 3024 6010 3080 6012
rect 3104 6010 3160 6012
rect 3184 6010 3240 6012
rect 3264 6010 3320 6012
rect 3024 5958 3070 6010
rect 3070 5958 3080 6010
rect 3104 5958 3134 6010
rect 3134 5958 3146 6010
rect 3146 5958 3160 6010
rect 3184 5958 3198 6010
rect 3198 5958 3210 6010
rect 3210 5958 3240 6010
rect 3264 5958 3274 6010
rect 3274 5958 3320 6010
rect 3024 5956 3080 5958
rect 3104 5956 3160 5958
rect 3184 5956 3240 5958
rect 3264 5956 3320 5958
rect 1950 5516 1952 5536
rect 1952 5516 2004 5536
rect 2004 5516 2006 5536
rect 1950 5480 2006 5516
rect 2305 5466 2361 5468
rect 2385 5466 2441 5468
rect 2465 5466 2521 5468
rect 2545 5466 2601 5468
rect 2305 5414 2351 5466
rect 2351 5414 2361 5466
rect 2385 5414 2415 5466
rect 2415 5414 2427 5466
rect 2427 5414 2441 5466
rect 2465 5414 2479 5466
rect 2479 5414 2491 5466
rect 2491 5414 2521 5466
rect 2545 5414 2555 5466
rect 2555 5414 2601 5466
rect 2305 5412 2361 5414
rect 2385 5412 2441 5414
rect 2465 5412 2521 5414
rect 2545 5412 2601 5414
rect 3684 5466 3740 5468
rect 3764 5466 3820 5468
rect 3844 5466 3900 5468
rect 3924 5466 3980 5468
rect 3684 5414 3730 5466
rect 3730 5414 3740 5466
rect 3764 5414 3794 5466
rect 3794 5414 3806 5466
rect 3806 5414 3820 5466
rect 3844 5414 3858 5466
rect 3858 5414 3870 5466
rect 3870 5414 3900 5466
rect 3924 5414 3934 5466
rect 3934 5414 3980 5466
rect 3684 5412 3740 5414
rect 3764 5412 3820 5414
rect 3844 5412 3900 5414
rect 3924 5412 3980 5414
rect 1645 4922 1701 4924
rect 1725 4922 1781 4924
rect 1805 4922 1861 4924
rect 1885 4922 1941 4924
rect 1645 4870 1691 4922
rect 1691 4870 1701 4922
rect 1725 4870 1755 4922
rect 1755 4870 1767 4922
rect 1767 4870 1781 4922
rect 1805 4870 1819 4922
rect 1819 4870 1831 4922
rect 1831 4870 1861 4922
rect 1885 4870 1895 4922
rect 1895 4870 1941 4922
rect 1645 4868 1701 4870
rect 1725 4868 1781 4870
rect 1805 4868 1861 4870
rect 1885 4868 1941 4870
rect 3024 4922 3080 4924
rect 3104 4922 3160 4924
rect 3184 4922 3240 4924
rect 3264 4922 3320 4924
rect 3024 4870 3070 4922
rect 3070 4870 3080 4922
rect 3104 4870 3134 4922
rect 3134 4870 3146 4922
rect 3146 4870 3160 4922
rect 3184 4870 3198 4922
rect 3198 4870 3210 4922
rect 3210 4870 3240 4922
rect 3264 4870 3274 4922
rect 3274 4870 3320 4922
rect 3024 4868 3080 4870
rect 3104 4868 3160 4870
rect 3184 4868 3240 4870
rect 3264 4868 3320 4870
rect 2305 4378 2361 4380
rect 2385 4378 2441 4380
rect 2465 4378 2521 4380
rect 2545 4378 2601 4380
rect 2305 4326 2351 4378
rect 2351 4326 2361 4378
rect 2385 4326 2415 4378
rect 2415 4326 2427 4378
rect 2427 4326 2441 4378
rect 2465 4326 2479 4378
rect 2479 4326 2491 4378
rect 2491 4326 2521 4378
rect 2545 4326 2555 4378
rect 2555 4326 2601 4378
rect 2305 4324 2361 4326
rect 2385 4324 2441 4326
rect 2465 4324 2521 4326
rect 2545 4324 2601 4326
rect 3684 4378 3740 4380
rect 3764 4378 3820 4380
rect 3844 4378 3900 4380
rect 3924 4378 3980 4380
rect 3684 4326 3730 4378
rect 3730 4326 3740 4378
rect 3764 4326 3794 4378
rect 3794 4326 3806 4378
rect 3806 4326 3820 4378
rect 3844 4326 3858 4378
rect 3858 4326 3870 4378
rect 3870 4326 3900 4378
rect 3924 4326 3934 4378
rect 3934 4326 3980 4378
rect 3684 4324 3740 4326
rect 3764 4324 3820 4326
rect 3844 4324 3900 4326
rect 3924 4324 3980 4326
rect 1645 3834 1701 3836
rect 1725 3834 1781 3836
rect 1805 3834 1861 3836
rect 1885 3834 1941 3836
rect 1645 3782 1691 3834
rect 1691 3782 1701 3834
rect 1725 3782 1755 3834
rect 1755 3782 1767 3834
rect 1767 3782 1781 3834
rect 1805 3782 1819 3834
rect 1819 3782 1831 3834
rect 1831 3782 1861 3834
rect 1885 3782 1895 3834
rect 1895 3782 1941 3834
rect 1645 3780 1701 3782
rect 1725 3780 1781 3782
rect 1805 3780 1861 3782
rect 1885 3780 1941 3782
rect 2305 3290 2361 3292
rect 2385 3290 2441 3292
rect 2465 3290 2521 3292
rect 2545 3290 2601 3292
rect 2305 3238 2351 3290
rect 2351 3238 2361 3290
rect 2385 3238 2415 3290
rect 2415 3238 2427 3290
rect 2427 3238 2441 3290
rect 2465 3238 2479 3290
rect 2479 3238 2491 3290
rect 2491 3238 2521 3290
rect 2545 3238 2555 3290
rect 2555 3238 2601 3290
rect 2305 3236 2361 3238
rect 2385 3236 2441 3238
rect 2465 3236 2521 3238
rect 2545 3236 2601 3238
rect 1645 2746 1701 2748
rect 1725 2746 1781 2748
rect 1805 2746 1861 2748
rect 1885 2746 1941 2748
rect 1645 2694 1691 2746
rect 1691 2694 1701 2746
rect 1725 2694 1755 2746
rect 1755 2694 1767 2746
rect 1767 2694 1781 2746
rect 1805 2694 1819 2746
rect 1819 2694 1831 2746
rect 1831 2694 1861 2746
rect 1885 2694 1895 2746
rect 1895 2694 1941 2746
rect 1645 2692 1701 2694
rect 1725 2692 1781 2694
rect 1805 2692 1861 2694
rect 1885 2692 1941 2694
rect 3024 3834 3080 3836
rect 3104 3834 3160 3836
rect 3184 3834 3240 3836
rect 3264 3834 3320 3836
rect 3024 3782 3070 3834
rect 3070 3782 3080 3834
rect 3104 3782 3134 3834
rect 3134 3782 3146 3834
rect 3146 3782 3160 3834
rect 3184 3782 3198 3834
rect 3198 3782 3210 3834
rect 3210 3782 3240 3834
rect 3264 3782 3274 3834
rect 3274 3782 3320 3834
rect 3024 3780 3080 3782
rect 3104 3780 3160 3782
rect 3184 3780 3240 3782
rect 3264 3780 3320 3782
rect 4403 6010 4459 6012
rect 4483 6010 4539 6012
rect 4563 6010 4619 6012
rect 4643 6010 4699 6012
rect 4403 5958 4449 6010
rect 4449 5958 4459 6010
rect 4483 5958 4513 6010
rect 4513 5958 4525 6010
rect 4525 5958 4539 6010
rect 4563 5958 4577 6010
rect 4577 5958 4589 6010
rect 4589 5958 4619 6010
rect 4643 5958 4653 6010
rect 4653 5958 4699 6010
rect 4403 5956 4459 5958
rect 4483 5956 4539 5958
rect 4563 5956 4619 5958
rect 4643 5956 4699 5958
rect 5782 6010 5838 6012
rect 5862 6010 5918 6012
rect 5942 6010 5998 6012
rect 6022 6010 6078 6012
rect 5782 5958 5828 6010
rect 5828 5958 5838 6010
rect 5862 5958 5892 6010
rect 5892 5958 5904 6010
rect 5904 5958 5918 6010
rect 5942 5958 5956 6010
rect 5956 5958 5968 6010
rect 5968 5958 5998 6010
rect 6022 5958 6032 6010
rect 6032 5958 6078 6010
rect 5782 5956 5838 5958
rect 5862 5956 5918 5958
rect 5942 5956 5998 5958
rect 6022 5956 6078 5958
rect 6274 5752 6330 5808
rect 5063 5466 5119 5468
rect 5143 5466 5199 5468
rect 5223 5466 5279 5468
rect 5303 5466 5359 5468
rect 5063 5414 5109 5466
rect 5109 5414 5119 5466
rect 5143 5414 5173 5466
rect 5173 5414 5185 5466
rect 5185 5414 5199 5466
rect 5223 5414 5237 5466
rect 5237 5414 5249 5466
rect 5249 5414 5279 5466
rect 5303 5414 5313 5466
rect 5313 5414 5359 5466
rect 5063 5412 5119 5414
rect 5143 5412 5199 5414
rect 5223 5412 5279 5414
rect 5303 5412 5359 5414
rect 6442 5466 6498 5468
rect 6522 5466 6578 5468
rect 6602 5466 6658 5468
rect 6682 5466 6738 5468
rect 6442 5414 6488 5466
rect 6488 5414 6498 5466
rect 6522 5414 6552 5466
rect 6552 5414 6564 5466
rect 6564 5414 6578 5466
rect 6602 5414 6616 5466
rect 6616 5414 6628 5466
rect 6628 5414 6658 5466
rect 6682 5414 6692 5466
rect 6692 5414 6738 5466
rect 6442 5412 6498 5414
rect 6522 5412 6578 5414
rect 6602 5412 6658 5414
rect 6682 5412 6738 5414
rect 4403 4922 4459 4924
rect 4483 4922 4539 4924
rect 4563 4922 4619 4924
rect 4643 4922 4699 4924
rect 4403 4870 4449 4922
rect 4449 4870 4459 4922
rect 4483 4870 4513 4922
rect 4513 4870 4525 4922
rect 4525 4870 4539 4922
rect 4563 4870 4577 4922
rect 4577 4870 4589 4922
rect 4589 4870 4619 4922
rect 4643 4870 4653 4922
rect 4653 4870 4699 4922
rect 4403 4868 4459 4870
rect 4483 4868 4539 4870
rect 4563 4868 4619 4870
rect 4643 4868 4699 4870
rect 4403 3834 4459 3836
rect 4483 3834 4539 3836
rect 4563 3834 4619 3836
rect 4643 3834 4699 3836
rect 4403 3782 4449 3834
rect 4449 3782 4459 3834
rect 4483 3782 4513 3834
rect 4513 3782 4525 3834
rect 4525 3782 4539 3834
rect 4563 3782 4577 3834
rect 4577 3782 4589 3834
rect 4589 3782 4619 3834
rect 4643 3782 4653 3834
rect 4653 3782 4699 3834
rect 4403 3780 4459 3782
rect 4483 3780 4539 3782
rect 4563 3780 4619 3782
rect 4643 3780 4699 3782
rect 3024 2746 3080 2748
rect 3104 2746 3160 2748
rect 3184 2746 3240 2748
rect 3264 2746 3320 2748
rect 3024 2694 3070 2746
rect 3070 2694 3080 2746
rect 3104 2694 3134 2746
rect 3134 2694 3146 2746
rect 3146 2694 3160 2746
rect 3184 2694 3198 2746
rect 3198 2694 3210 2746
rect 3210 2694 3240 2746
rect 3264 2694 3274 2746
rect 3274 2694 3320 2746
rect 3024 2692 3080 2694
rect 3104 2692 3160 2694
rect 3184 2692 3240 2694
rect 3264 2692 3320 2694
rect 3684 3290 3740 3292
rect 3764 3290 3820 3292
rect 3844 3290 3900 3292
rect 3924 3290 3980 3292
rect 3684 3238 3730 3290
rect 3730 3238 3740 3290
rect 3764 3238 3794 3290
rect 3794 3238 3806 3290
rect 3806 3238 3820 3290
rect 3844 3238 3858 3290
rect 3858 3238 3870 3290
rect 3870 3238 3900 3290
rect 3924 3238 3934 3290
rect 3934 3238 3980 3290
rect 3684 3236 3740 3238
rect 3764 3236 3820 3238
rect 3844 3236 3900 3238
rect 3924 3236 3980 3238
rect 5782 4922 5838 4924
rect 5862 4922 5918 4924
rect 5942 4922 5998 4924
rect 6022 4922 6078 4924
rect 5782 4870 5828 4922
rect 5828 4870 5838 4922
rect 5862 4870 5892 4922
rect 5892 4870 5904 4922
rect 5904 4870 5918 4922
rect 5942 4870 5956 4922
rect 5956 4870 5968 4922
rect 5968 4870 5998 4922
rect 6022 4870 6032 4922
rect 6032 4870 6078 4922
rect 5782 4868 5838 4870
rect 5862 4868 5918 4870
rect 5942 4868 5998 4870
rect 6022 4868 6078 4870
rect 6182 4800 6238 4856
rect 5063 4378 5119 4380
rect 5143 4378 5199 4380
rect 5223 4378 5279 4380
rect 5303 4378 5359 4380
rect 5063 4326 5109 4378
rect 5109 4326 5119 4378
rect 5143 4326 5173 4378
rect 5173 4326 5185 4378
rect 5185 4326 5199 4378
rect 5223 4326 5237 4378
rect 5237 4326 5249 4378
rect 5249 4326 5279 4378
rect 5303 4326 5313 4378
rect 5313 4326 5359 4378
rect 5063 4324 5119 4326
rect 5143 4324 5199 4326
rect 5223 4324 5279 4326
rect 5303 4324 5359 4326
rect 6442 4378 6498 4380
rect 6522 4378 6578 4380
rect 6602 4378 6658 4380
rect 6682 4378 6738 4380
rect 6442 4326 6488 4378
rect 6488 4326 6498 4378
rect 6522 4326 6552 4378
rect 6552 4326 6564 4378
rect 6564 4326 6578 4378
rect 6602 4326 6616 4378
rect 6616 4326 6628 4378
rect 6628 4326 6658 4378
rect 6682 4326 6692 4378
rect 6692 4326 6738 4378
rect 6442 4324 6498 4326
rect 6522 4324 6578 4326
rect 6602 4324 6658 4326
rect 6682 4324 6738 4326
rect 6274 4120 6330 4176
rect 5782 3834 5838 3836
rect 5862 3834 5918 3836
rect 5942 3834 5998 3836
rect 6022 3834 6078 3836
rect 5782 3782 5828 3834
rect 5828 3782 5838 3834
rect 5862 3782 5892 3834
rect 5892 3782 5904 3834
rect 5904 3782 5918 3834
rect 5942 3782 5956 3834
rect 5956 3782 5968 3834
rect 5968 3782 5998 3834
rect 6022 3782 6032 3834
rect 6032 3782 6078 3834
rect 5782 3780 5838 3782
rect 5862 3780 5918 3782
rect 5942 3780 5998 3782
rect 6022 3780 6078 3782
rect 6182 3440 6238 3496
rect 5063 3290 5119 3292
rect 5143 3290 5199 3292
rect 5223 3290 5279 3292
rect 5303 3290 5359 3292
rect 5063 3238 5109 3290
rect 5109 3238 5119 3290
rect 5143 3238 5173 3290
rect 5173 3238 5185 3290
rect 5185 3238 5199 3290
rect 5223 3238 5237 3290
rect 5237 3238 5249 3290
rect 5249 3238 5279 3290
rect 5303 3238 5313 3290
rect 5313 3238 5359 3290
rect 5063 3236 5119 3238
rect 5143 3236 5199 3238
rect 5223 3236 5279 3238
rect 5303 3236 5359 3238
rect 6442 3290 6498 3292
rect 6522 3290 6578 3292
rect 6602 3290 6658 3292
rect 6682 3290 6738 3292
rect 6442 3238 6488 3290
rect 6488 3238 6498 3290
rect 6522 3238 6552 3290
rect 6552 3238 6564 3290
rect 6564 3238 6578 3290
rect 6602 3238 6616 3290
rect 6616 3238 6628 3290
rect 6628 3238 6658 3290
rect 6682 3238 6692 3290
rect 6692 3238 6738 3290
rect 6442 3236 6498 3238
rect 6522 3236 6578 3238
rect 6602 3236 6658 3238
rect 6682 3236 6738 3238
rect 4403 2746 4459 2748
rect 4483 2746 4539 2748
rect 4563 2746 4619 2748
rect 4643 2746 4699 2748
rect 4403 2694 4449 2746
rect 4449 2694 4459 2746
rect 4483 2694 4513 2746
rect 4513 2694 4525 2746
rect 4525 2694 4539 2746
rect 4563 2694 4577 2746
rect 4577 2694 4589 2746
rect 4589 2694 4619 2746
rect 4643 2694 4653 2746
rect 4653 2694 4699 2746
rect 4403 2692 4459 2694
rect 4483 2692 4539 2694
rect 4563 2692 4619 2694
rect 4643 2692 4699 2694
rect 5782 2746 5838 2748
rect 5862 2746 5918 2748
rect 5942 2746 5998 2748
rect 6022 2746 6078 2748
rect 5782 2694 5828 2746
rect 5828 2694 5838 2746
rect 5862 2694 5892 2746
rect 5892 2694 5904 2746
rect 5904 2694 5918 2746
rect 5942 2694 5956 2746
rect 5956 2694 5968 2746
rect 5968 2694 5998 2746
rect 6022 2694 6032 2746
rect 6032 2694 6078 2746
rect 5782 2692 5838 2694
rect 5862 2692 5918 2694
rect 5942 2692 5998 2694
rect 6022 2692 6078 2694
rect 2305 2202 2361 2204
rect 2385 2202 2441 2204
rect 2465 2202 2521 2204
rect 2545 2202 2601 2204
rect 2305 2150 2351 2202
rect 2351 2150 2361 2202
rect 2385 2150 2415 2202
rect 2415 2150 2427 2202
rect 2427 2150 2441 2202
rect 2465 2150 2479 2202
rect 2479 2150 2491 2202
rect 2491 2150 2521 2202
rect 2545 2150 2555 2202
rect 2555 2150 2601 2202
rect 2305 2148 2361 2150
rect 2385 2148 2441 2150
rect 2465 2148 2521 2150
rect 2545 2148 2601 2150
rect 3684 2202 3740 2204
rect 3764 2202 3820 2204
rect 3844 2202 3900 2204
rect 3924 2202 3980 2204
rect 3684 2150 3730 2202
rect 3730 2150 3740 2202
rect 3764 2150 3794 2202
rect 3794 2150 3806 2202
rect 3806 2150 3820 2202
rect 3844 2150 3858 2202
rect 3858 2150 3870 2202
rect 3870 2150 3900 2202
rect 3924 2150 3934 2202
rect 3934 2150 3980 2202
rect 3684 2148 3740 2150
rect 3764 2148 3820 2150
rect 3844 2148 3900 2150
rect 3924 2148 3980 2150
rect 5063 2202 5119 2204
rect 5143 2202 5199 2204
rect 5223 2202 5279 2204
rect 5303 2202 5359 2204
rect 5063 2150 5109 2202
rect 5109 2150 5119 2202
rect 5143 2150 5173 2202
rect 5173 2150 5185 2202
rect 5185 2150 5199 2202
rect 5223 2150 5237 2202
rect 5237 2150 5249 2202
rect 5249 2150 5279 2202
rect 5303 2150 5313 2202
rect 5313 2150 5359 2202
rect 5063 2148 5119 2150
rect 5143 2148 5199 2150
rect 5223 2148 5279 2150
rect 5303 2148 5359 2150
rect 6442 2202 6498 2204
rect 6522 2202 6578 2204
rect 6602 2202 6658 2204
rect 6682 2202 6738 2204
rect 6442 2150 6488 2202
rect 6488 2150 6498 2202
rect 6522 2150 6552 2202
rect 6552 2150 6564 2202
rect 6564 2150 6578 2202
rect 6602 2150 6616 2202
rect 6616 2150 6628 2202
rect 6628 2150 6658 2202
rect 6682 2150 6692 2202
rect 6692 2150 6738 2202
rect 6442 2148 6498 2150
rect 6522 2148 6578 2150
rect 6602 2148 6658 2150
rect 6682 2148 6738 2150
<< metal3 >>
rect 2295 7648 2611 7649
rect 0 7578 800 7608
rect 2295 7584 2301 7648
rect 2365 7584 2381 7648
rect 2445 7584 2461 7648
rect 2525 7584 2541 7648
rect 2605 7584 2611 7648
rect 2295 7583 2611 7584
rect 3674 7648 3990 7649
rect 3674 7584 3680 7648
rect 3744 7584 3760 7648
rect 3824 7584 3840 7648
rect 3904 7584 3920 7648
rect 3984 7584 3990 7648
rect 3674 7583 3990 7584
rect 5053 7648 5369 7649
rect 5053 7584 5059 7648
rect 5123 7584 5139 7648
rect 5203 7584 5219 7648
rect 5283 7584 5299 7648
rect 5363 7584 5369 7648
rect 5053 7583 5369 7584
rect 6432 7648 6748 7649
rect 6432 7584 6438 7648
rect 6502 7584 6518 7648
rect 6582 7584 6598 7648
rect 6662 7584 6678 7648
rect 6742 7584 6748 7648
rect 6432 7583 6748 7584
rect 0 7488 858 7578
rect 798 7445 858 7488
rect 798 7440 907 7445
rect 798 7384 846 7440
rect 902 7384 907 7440
rect 798 7382 907 7384
rect 841 7379 907 7382
rect 1635 7104 1951 7105
rect 1635 7040 1641 7104
rect 1705 7040 1721 7104
rect 1785 7040 1801 7104
rect 1865 7040 1881 7104
rect 1945 7040 1951 7104
rect 1635 7039 1951 7040
rect 3014 7104 3330 7105
rect 3014 7040 3020 7104
rect 3084 7040 3100 7104
rect 3164 7040 3180 7104
rect 3244 7040 3260 7104
rect 3324 7040 3330 7104
rect 3014 7039 3330 7040
rect 4393 7104 4709 7105
rect 4393 7040 4399 7104
rect 4463 7040 4479 7104
rect 4543 7040 4559 7104
rect 4623 7040 4639 7104
rect 4703 7040 4709 7104
rect 4393 7039 4709 7040
rect 5772 7104 6088 7105
rect 5772 7040 5778 7104
rect 5842 7040 5858 7104
rect 5922 7040 5938 7104
rect 6002 7040 6018 7104
rect 6082 7040 6088 7104
rect 5772 7039 6088 7040
rect 0 6898 800 6928
rect 1485 6898 1551 6901
rect 0 6896 1551 6898
rect 0 6840 1490 6896
rect 1546 6840 1551 6896
rect 0 6838 1551 6840
rect 0 6808 800 6838
rect 1485 6835 1551 6838
rect 2295 6560 2611 6561
rect 2295 6496 2301 6560
rect 2365 6496 2381 6560
rect 2445 6496 2461 6560
rect 2525 6496 2541 6560
rect 2605 6496 2611 6560
rect 2295 6495 2611 6496
rect 3674 6560 3990 6561
rect 3674 6496 3680 6560
rect 3744 6496 3760 6560
rect 3824 6496 3840 6560
rect 3904 6496 3920 6560
rect 3984 6496 3990 6560
rect 3674 6495 3990 6496
rect 5053 6560 5369 6561
rect 5053 6496 5059 6560
rect 5123 6496 5139 6560
rect 5203 6496 5219 6560
rect 5283 6496 5299 6560
rect 5363 6496 5369 6560
rect 5053 6495 5369 6496
rect 6432 6560 6748 6561
rect 6432 6496 6438 6560
rect 6502 6496 6518 6560
rect 6582 6496 6598 6560
rect 6662 6496 6678 6560
rect 6742 6496 6748 6560
rect 6432 6495 6748 6496
rect 0 6218 800 6248
rect 1209 6218 1275 6221
rect 0 6216 1275 6218
rect 0 6160 1214 6216
rect 1270 6160 1275 6216
rect 0 6158 1275 6160
rect 0 6128 800 6158
rect 1209 6155 1275 6158
rect 1635 6016 1951 6017
rect 1635 5952 1641 6016
rect 1705 5952 1721 6016
rect 1785 5952 1801 6016
rect 1865 5952 1881 6016
rect 1945 5952 1951 6016
rect 1635 5951 1951 5952
rect 3014 6016 3330 6017
rect 3014 5952 3020 6016
rect 3084 5952 3100 6016
rect 3164 5952 3180 6016
rect 3244 5952 3260 6016
rect 3324 5952 3330 6016
rect 3014 5951 3330 5952
rect 4393 6016 4709 6017
rect 4393 5952 4399 6016
rect 4463 5952 4479 6016
rect 4543 5952 4559 6016
rect 4623 5952 4639 6016
rect 4703 5952 4709 6016
rect 4393 5951 4709 5952
rect 5772 6016 6088 6017
rect 5772 5952 5778 6016
rect 5842 5952 5858 6016
rect 5922 5952 5938 6016
rect 6002 5952 6018 6016
rect 6082 5952 6088 6016
rect 5772 5951 6088 5952
rect 6269 5810 6335 5813
rect 6862 5810 6868 5812
rect 6269 5808 6868 5810
rect 6269 5752 6274 5808
rect 6330 5752 6868 5808
rect 6269 5750 6868 5752
rect 6269 5747 6335 5750
rect 6862 5748 6868 5750
rect 6932 5748 6938 5812
rect 0 5538 800 5568
rect 1945 5538 2011 5541
rect 6933 5540 7733 5568
rect 0 5536 2011 5538
rect 0 5480 1950 5536
rect 2006 5480 2011 5536
rect 0 5478 2011 5480
rect 0 5448 800 5478
rect 1945 5475 2011 5478
rect 6862 5476 6868 5540
rect 6932 5476 7733 5540
rect 2295 5472 2611 5473
rect 2295 5408 2301 5472
rect 2365 5408 2381 5472
rect 2445 5408 2461 5472
rect 2525 5408 2541 5472
rect 2605 5408 2611 5472
rect 2295 5407 2611 5408
rect 3674 5472 3990 5473
rect 3674 5408 3680 5472
rect 3744 5408 3760 5472
rect 3824 5408 3840 5472
rect 3904 5408 3920 5472
rect 3984 5408 3990 5472
rect 3674 5407 3990 5408
rect 5053 5472 5369 5473
rect 5053 5408 5059 5472
rect 5123 5408 5139 5472
rect 5203 5408 5219 5472
rect 5283 5408 5299 5472
rect 5363 5408 5369 5472
rect 5053 5407 5369 5408
rect 6432 5472 6748 5473
rect 6432 5408 6438 5472
rect 6502 5408 6518 5472
rect 6582 5408 6598 5472
rect 6662 5408 6678 5472
rect 6742 5408 6748 5472
rect 6933 5448 7733 5476
rect 6432 5407 6748 5408
rect 1635 4928 1951 4929
rect 1635 4864 1641 4928
rect 1705 4864 1721 4928
rect 1785 4864 1801 4928
rect 1865 4864 1881 4928
rect 1945 4864 1951 4928
rect 1635 4863 1951 4864
rect 3014 4928 3330 4929
rect 3014 4864 3020 4928
rect 3084 4864 3100 4928
rect 3164 4864 3180 4928
rect 3244 4864 3260 4928
rect 3324 4864 3330 4928
rect 3014 4863 3330 4864
rect 4393 4928 4709 4929
rect 4393 4864 4399 4928
rect 4463 4864 4479 4928
rect 4543 4864 4559 4928
rect 4623 4864 4639 4928
rect 4703 4864 4709 4928
rect 4393 4863 4709 4864
rect 5772 4928 6088 4929
rect 5772 4864 5778 4928
rect 5842 4864 5858 4928
rect 5922 4864 5938 4928
rect 6002 4864 6018 4928
rect 6082 4864 6088 4928
rect 5772 4863 6088 4864
rect 6177 4858 6243 4861
rect 6933 4858 7733 4888
rect 6177 4856 7733 4858
rect 6177 4800 6182 4856
rect 6238 4800 7733 4856
rect 6177 4798 7733 4800
rect 6177 4795 6243 4798
rect 6933 4768 7733 4798
rect 2295 4384 2611 4385
rect 2295 4320 2301 4384
rect 2365 4320 2381 4384
rect 2445 4320 2461 4384
rect 2525 4320 2541 4384
rect 2605 4320 2611 4384
rect 2295 4319 2611 4320
rect 3674 4384 3990 4385
rect 3674 4320 3680 4384
rect 3744 4320 3760 4384
rect 3824 4320 3840 4384
rect 3904 4320 3920 4384
rect 3984 4320 3990 4384
rect 3674 4319 3990 4320
rect 5053 4384 5369 4385
rect 5053 4320 5059 4384
rect 5123 4320 5139 4384
rect 5203 4320 5219 4384
rect 5283 4320 5299 4384
rect 5363 4320 5369 4384
rect 5053 4319 5369 4320
rect 6432 4384 6748 4385
rect 6432 4320 6438 4384
rect 6502 4320 6518 4384
rect 6582 4320 6598 4384
rect 6662 4320 6678 4384
rect 6742 4320 6748 4384
rect 6432 4319 6748 4320
rect 6269 4178 6335 4181
rect 6933 4178 7733 4208
rect 6269 4176 7733 4178
rect 6269 4120 6274 4176
rect 6330 4120 7733 4176
rect 6269 4118 7733 4120
rect 6269 4115 6335 4118
rect 6933 4088 7733 4118
rect 1635 3840 1951 3841
rect 1635 3776 1641 3840
rect 1705 3776 1721 3840
rect 1785 3776 1801 3840
rect 1865 3776 1881 3840
rect 1945 3776 1951 3840
rect 1635 3775 1951 3776
rect 3014 3840 3330 3841
rect 3014 3776 3020 3840
rect 3084 3776 3100 3840
rect 3164 3776 3180 3840
rect 3244 3776 3260 3840
rect 3324 3776 3330 3840
rect 3014 3775 3330 3776
rect 4393 3840 4709 3841
rect 4393 3776 4399 3840
rect 4463 3776 4479 3840
rect 4543 3776 4559 3840
rect 4623 3776 4639 3840
rect 4703 3776 4709 3840
rect 4393 3775 4709 3776
rect 5772 3840 6088 3841
rect 5772 3776 5778 3840
rect 5842 3776 5858 3840
rect 5922 3776 5938 3840
rect 6002 3776 6018 3840
rect 6082 3776 6088 3840
rect 5772 3775 6088 3776
rect 6177 3498 6243 3501
rect 6933 3498 7733 3528
rect 6177 3496 7733 3498
rect 6177 3440 6182 3496
rect 6238 3440 7733 3496
rect 6177 3438 7733 3440
rect 6177 3435 6243 3438
rect 6933 3408 7733 3438
rect 2295 3296 2611 3297
rect 2295 3232 2301 3296
rect 2365 3232 2381 3296
rect 2445 3232 2461 3296
rect 2525 3232 2541 3296
rect 2605 3232 2611 3296
rect 2295 3231 2611 3232
rect 3674 3296 3990 3297
rect 3674 3232 3680 3296
rect 3744 3232 3760 3296
rect 3824 3232 3840 3296
rect 3904 3232 3920 3296
rect 3984 3232 3990 3296
rect 3674 3231 3990 3232
rect 5053 3296 5369 3297
rect 5053 3232 5059 3296
rect 5123 3232 5139 3296
rect 5203 3232 5219 3296
rect 5283 3232 5299 3296
rect 5363 3232 5369 3296
rect 5053 3231 5369 3232
rect 6432 3296 6748 3297
rect 6432 3232 6438 3296
rect 6502 3232 6518 3296
rect 6582 3232 6598 3296
rect 6662 3232 6678 3296
rect 6742 3232 6748 3296
rect 6432 3231 6748 3232
rect 1635 2752 1951 2753
rect 1635 2688 1641 2752
rect 1705 2688 1721 2752
rect 1785 2688 1801 2752
rect 1865 2688 1881 2752
rect 1945 2688 1951 2752
rect 1635 2687 1951 2688
rect 3014 2752 3330 2753
rect 3014 2688 3020 2752
rect 3084 2688 3100 2752
rect 3164 2688 3180 2752
rect 3244 2688 3260 2752
rect 3324 2688 3330 2752
rect 3014 2687 3330 2688
rect 4393 2752 4709 2753
rect 4393 2688 4399 2752
rect 4463 2688 4479 2752
rect 4543 2688 4559 2752
rect 4623 2688 4639 2752
rect 4703 2688 4709 2752
rect 4393 2687 4709 2688
rect 5772 2752 6088 2753
rect 5772 2688 5778 2752
rect 5842 2688 5858 2752
rect 5922 2688 5938 2752
rect 6002 2688 6018 2752
rect 6082 2688 6088 2752
rect 5772 2687 6088 2688
rect 2295 2208 2611 2209
rect 2295 2144 2301 2208
rect 2365 2144 2381 2208
rect 2445 2144 2461 2208
rect 2525 2144 2541 2208
rect 2605 2144 2611 2208
rect 2295 2143 2611 2144
rect 3674 2208 3990 2209
rect 3674 2144 3680 2208
rect 3744 2144 3760 2208
rect 3824 2144 3840 2208
rect 3904 2144 3920 2208
rect 3984 2144 3990 2208
rect 3674 2143 3990 2144
rect 5053 2208 5369 2209
rect 5053 2144 5059 2208
rect 5123 2144 5139 2208
rect 5203 2144 5219 2208
rect 5283 2144 5299 2208
rect 5363 2144 5369 2208
rect 5053 2143 5369 2144
rect 6432 2208 6748 2209
rect 6432 2144 6438 2208
rect 6502 2144 6518 2208
rect 6582 2144 6598 2208
rect 6662 2144 6678 2208
rect 6742 2144 6748 2208
rect 6432 2143 6748 2144
<< via3 >>
rect 2301 7644 2365 7648
rect 2301 7588 2305 7644
rect 2305 7588 2361 7644
rect 2361 7588 2365 7644
rect 2301 7584 2365 7588
rect 2381 7644 2445 7648
rect 2381 7588 2385 7644
rect 2385 7588 2441 7644
rect 2441 7588 2445 7644
rect 2381 7584 2445 7588
rect 2461 7644 2525 7648
rect 2461 7588 2465 7644
rect 2465 7588 2521 7644
rect 2521 7588 2525 7644
rect 2461 7584 2525 7588
rect 2541 7644 2605 7648
rect 2541 7588 2545 7644
rect 2545 7588 2601 7644
rect 2601 7588 2605 7644
rect 2541 7584 2605 7588
rect 3680 7644 3744 7648
rect 3680 7588 3684 7644
rect 3684 7588 3740 7644
rect 3740 7588 3744 7644
rect 3680 7584 3744 7588
rect 3760 7644 3824 7648
rect 3760 7588 3764 7644
rect 3764 7588 3820 7644
rect 3820 7588 3824 7644
rect 3760 7584 3824 7588
rect 3840 7644 3904 7648
rect 3840 7588 3844 7644
rect 3844 7588 3900 7644
rect 3900 7588 3904 7644
rect 3840 7584 3904 7588
rect 3920 7644 3984 7648
rect 3920 7588 3924 7644
rect 3924 7588 3980 7644
rect 3980 7588 3984 7644
rect 3920 7584 3984 7588
rect 5059 7644 5123 7648
rect 5059 7588 5063 7644
rect 5063 7588 5119 7644
rect 5119 7588 5123 7644
rect 5059 7584 5123 7588
rect 5139 7644 5203 7648
rect 5139 7588 5143 7644
rect 5143 7588 5199 7644
rect 5199 7588 5203 7644
rect 5139 7584 5203 7588
rect 5219 7644 5283 7648
rect 5219 7588 5223 7644
rect 5223 7588 5279 7644
rect 5279 7588 5283 7644
rect 5219 7584 5283 7588
rect 5299 7644 5363 7648
rect 5299 7588 5303 7644
rect 5303 7588 5359 7644
rect 5359 7588 5363 7644
rect 5299 7584 5363 7588
rect 6438 7644 6502 7648
rect 6438 7588 6442 7644
rect 6442 7588 6498 7644
rect 6498 7588 6502 7644
rect 6438 7584 6502 7588
rect 6518 7644 6582 7648
rect 6518 7588 6522 7644
rect 6522 7588 6578 7644
rect 6578 7588 6582 7644
rect 6518 7584 6582 7588
rect 6598 7644 6662 7648
rect 6598 7588 6602 7644
rect 6602 7588 6658 7644
rect 6658 7588 6662 7644
rect 6598 7584 6662 7588
rect 6678 7644 6742 7648
rect 6678 7588 6682 7644
rect 6682 7588 6738 7644
rect 6738 7588 6742 7644
rect 6678 7584 6742 7588
rect 1641 7100 1705 7104
rect 1641 7044 1645 7100
rect 1645 7044 1701 7100
rect 1701 7044 1705 7100
rect 1641 7040 1705 7044
rect 1721 7100 1785 7104
rect 1721 7044 1725 7100
rect 1725 7044 1781 7100
rect 1781 7044 1785 7100
rect 1721 7040 1785 7044
rect 1801 7100 1865 7104
rect 1801 7044 1805 7100
rect 1805 7044 1861 7100
rect 1861 7044 1865 7100
rect 1801 7040 1865 7044
rect 1881 7100 1945 7104
rect 1881 7044 1885 7100
rect 1885 7044 1941 7100
rect 1941 7044 1945 7100
rect 1881 7040 1945 7044
rect 3020 7100 3084 7104
rect 3020 7044 3024 7100
rect 3024 7044 3080 7100
rect 3080 7044 3084 7100
rect 3020 7040 3084 7044
rect 3100 7100 3164 7104
rect 3100 7044 3104 7100
rect 3104 7044 3160 7100
rect 3160 7044 3164 7100
rect 3100 7040 3164 7044
rect 3180 7100 3244 7104
rect 3180 7044 3184 7100
rect 3184 7044 3240 7100
rect 3240 7044 3244 7100
rect 3180 7040 3244 7044
rect 3260 7100 3324 7104
rect 3260 7044 3264 7100
rect 3264 7044 3320 7100
rect 3320 7044 3324 7100
rect 3260 7040 3324 7044
rect 4399 7100 4463 7104
rect 4399 7044 4403 7100
rect 4403 7044 4459 7100
rect 4459 7044 4463 7100
rect 4399 7040 4463 7044
rect 4479 7100 4543 7104
rect 4479 7044 4483 7100
rect 4483 7044 4539 7100
rect 4539 7044 4543 7100
rect 4479 7040 4543 7044
rect 4559 7100 4623 7104
rect 4559 7044 4563 7100
rect 4563 7044 4619 7100
rect 4619 7044 4623 7100
rect 4559 7040 4623 7044
rect 4639 7100 4703 7104
rect 4639 7044 4643 7100
rect 4643 7044 4699 7100
rect 4699 7044 4703 7100
rect 4639 7040 4703 7044
rect 5778 7100 5842 7104
rect 5778 7044 5782 7100
rect 5782 7044 5838 7100
rect 5838 7044 5842 7100
rect 5778 7040 5842 7044
rect 5858 7100 5922 7104
rect 5858 7044 5862 7100
rect 5862 7044 5918 7100
rect 5918 7044 5922 7100
rect 5858 7040 5922 7044
rect 5938 7100 6002 7104
rect 5938 7044 5942 7100
rect 5942 7044 5998 7100
rect 5998 7044 6002 7100
rect 5938 7040 6002 7044
rect 6018 7100 6082 7104
rect 6018 7044 6022 7100
rect 6022 7044 6078 7100
rect 6078 7044 6082 7100
rect 6018 7040 6082 7044
rect 2301 6556 2365 6560
rect 2301 6500 2305 6556
rect 2305 6500 2361 6556
rect 2361 6500 2365 6556
rect 2301 6496 2365 6500
rect 2381 6556 2445 6560
rect 2381 6500 2385 6556
rect 2385 6500 2441 6556
rect 2441 6500 2445 6556
rect 2381 6496 2445 6500
rect 2461 6556 2525 6560
rect 2461 6500 2465 6556
rect 2465 6500 2521 6556
rect 2521 6500 2525 6556
rect 2461 6496 2525 6500
rect 2541 6556 2605 6560
rect 2541 6500 2545 6556
rect 2545 6500 2601 6556
rect 2601 6500 2605 6556
rect 2541 6496 2605 6500
rect 3680 6556 3744 6560
rect 3680 6500 3684 6556
rect 3684 6500 3740 6556
rect 3740 6500 3744 6556
rect 3680 6496 3744 6500
rect 3760 6556 3824 6560
rect 3760 6500 3764 6556
rect 3764 6500 3820 6556
rect 3820 6500 3824 6556
rect 3760 6496 3824 6500
rect 3840 6556 3904 6560
rect 3840 6500 3844 6556
rect 3844 6500 3900 6556
rect 3900 6500 3904 6556
rect 3840 6496 3904 6500
rect 3920 6556 3984 6560
rect 3920 6500 3924 6556
rect 3924 6500 3980 6556
rect 3980 6500 3984 6556
rect 3920 6496 3984 6500
rect 5059 6556 5123 6560
rect 5059 6500 5063 6556
rect 5063 6500 5119 6556
rect 5119 6500 5123 6556
rect 5059 6496 5123 6500
rect 5139 6556 5203 6560
rect 5139 6500 5143 6556
rect 5143 6500 5199 6556
rect 5199 6500 5203 6556
rect 5139 6496 5203 6500
rect 5219 6556 5283 6560
rect 5219 6500 5223 6556
rect 5223 6500 5279 6556
rect 5279 6500 5283 6556
rect 5219 6496 5283 6500
rect 5299 6556 5363 6560
rect 5299 6500 5303 6556
rect 5303 6500 5359 6556
rect 5359 6500 5363 6556
rect 5299 6496 5363 6500
rect 6438 6556 6502 6560
rect 6438 6500 6442 6556
rect 6442 6500 6498 6556
rect 6498 6500 6502 6556
rect 6438 6496 6502 6500
rect 6518 6556 6582 6560
rect 6518 6500 6522 6556
rect 6522 6500 6578 6556
rect 6578 6500 6582 6556
rect 6518 6496 6582 6500
rect 6598 6556 6662 6560
rect 6598 6500 6602 6556
rect 6602 6500 6658 6556
rect 6658 6500 6662 6556
rect 6598 6496 6662 6500
rect 6678 6556 6742 6560
rect 6678 6500 6682 6556
rect 6682 6500 6738 6556
rect 6738 6500 6742 6556
rect 6678 6496 6742 6500
rect 1641 6012 1705 6016
rect 1641 5956 1645 6012
rect 1645 5956 1701 6012
rect 1701 5956 1705 6012
rect 1641 5952 1705 5956
rect 1721 6012 1785 6016
rect 1721 5956 1725 6012
rect 1725 5956 1781 6012
rect 1781 5956 1785 6012
rect 1721 5952 1785 5956
rect 1801 6012 1865 6016
rect 1801 5956 1805 6012
rect 1805 5956 1861 6012
rect 1861 5956 1865 6012
rect 1801 5952 1865 5956
rect 1881 6012 1945 6016
rect 1881 5956 1885 6012
rect 1885 5956 1941 6012
rect 1941 5956 1945 6012
rect 1881 5952 1945 5956
rect 3020 6012 3084 6016
rect 3020 5956 3024 6012
rect 3024 5956 3080 6012
rect 3080 5956 3084 6012
rect 3020 5952 3084 5956
rect 3100 6012 3164 6016
rect 3100 5956 3104 6012
rect 3104 5956 3160 6012
rect 3160 5956 3164 6012
rect 3100 5952 3164 5956
rect 3180 6012 3244 6016
rect 3180 5956 3184 6012
rect 3184 5956 3240 6012
rect 3240 5956 3244 6012
rect 3180 5952 3244 5956
rect 3260 6012 3324 6016
rect 3260 5956 3264 6012
rect 3264 5956 3320 6012
rect 3320 5956 3324 6012
rect 3260 5952 3324 5956
rect 4399 6012 4463 6016
rect 4399 5956 4403 6012
rect 4403 5956 4459 6012
rect 4459 5956 4463 6012
rect 4399 5952 4463 5956
rect 4479 6012 4543 6016
rect 4479 5956 4483 6012
rect 4483 5956 4539 6012
rect 4539 5956 4543 6012
rect 4479 5952 4543 5956
rect 4559 6012 4623 6016
rect 4559 5956 4563 6012
rect 4563 5956 4619 6012
rect 4619 5956 4623 6012
rect 4559 5952 4623 5956
rect 4639 6012 4703 6016
rect 4639 5956 4643 6012
rect 4643 5956 4699 6012
rect 4699 5956 4703 6012
rect 4639 5952 4703 5956
rect 5778 6012 5842 6016
rect 5778 5956 5782 6012
rect 5782 5956 5838 6012
rect 5838 5956 5842 6012
rect 5778 5952 5842 5956
rect 5858 6012 5922 6016
rect 5858 5956 5862 6012
rect 5862 5956 5918 6012
rect 5918 5956 5922 6012
rect 5858 5952 5922 5956
rect 5938 6012 6002 6016
rect 5938 5956 5942 6012
rect 5942 5956 5998 6012
rect 5998 5956 6002 6012
rect 5938 5952 6002 5956
rect 6018 6012 6082 6016
rect 6018 5956 6022 6012
rect 6022 5956 6078 6012
rect 6078 5956 6082 6012
rect 6018 5952 6082 5956
rect 6868 5748 6932 5812
rect 6868 5476 6932 5540
rect 2301 5468 2365 5472
rect 2301 5412 2305 5468
rect 2305 5412 2361 5468
rect 2361 5412 2365 5468
rect 2301 5408 2365 5412
rect 2381 5468 2445 5472
rect 2381 5412 2385 5468
rect 2385 5412 2441 5468
rect 2441 5412 2445 5468
rect 2381 5408 2445 5412
rect 2461 5468 2525 5472
rect 2461 5412 2465 5468
rect 2465 5412 2521 5468
rect 2521 5412 2525 5468
rect 2461 5408 2525 5412
rect 2541 5468 2605 5472
rect 2541 5412 2545 5468
rect 2545 5412 2601 5468
rect 2601 5412 2605 5468
rect 2541 5408 2605 5412
rect 3680 5468 3744 5472
rect 3680 5412 3684 5468
rect 3684 5412 3740 5468
rect 3740 5412 3744 5468
rect 3680 5408 3744 5412
rect 3760 5468 3824 5472
rect 3760 5412 3764 5468
rect 3764 5412 3820 5468
rect 3820 5412 3824 5468
rect 3760 5408 3824 5412
rect 3840 5468 3904 5472
rect 3840 5412 3844 5468
rect 3844 5412 3900 5468
rect 3900 5412 3904 5468
rect 3840 5408 3904 5412
rect 3920 5468 3984 5472
rect 3920 5412 3924 5468
rect 3924 5412 3980 5468
rect 3980 5412 3984 5468
rect 3920 5408 3984 5412
rect 5059 5468 5123 5472
rect 5059 5412 5063 5468
rect 5063 5412 5119 5468
rect 5119 5412 5123 5468
rect 5059 5408 5123 5412
rect 5139 5468 5203 5472
rect 5139 5412 5143 5468
rect 5143 5412 5199 5468
rect 5199 5412 5203 5468
rect 5139 5408 5203 5412
rect 5219 5468 5283 5472
rect 5219 5412 5223 5468
rect 5223 5412 5279 5468
rect 5279 5412 5283 5468
rect 5219 5408 5283 5412
rect 5299 5468 5363 5472
rect 5299 5412 5303 5468
rect 5303 5412 5359 5468
rect 5359 5412 5363 5468
rect 5299 5408 5363 5412
rect 6438 5468 6502 5472
rect 6438 5412 6442 5468
rect 6442 5412 6498 5468
rect 6498 5412 6502 5468
rect 6438 5408 6502 5412
rect 6518 5468 6582 5472
rect 6518 5412 6522 5468
rect 6522 5412 6578 5468
rect 6578 5412 6582 5468
rect 6518 5408 6582 5412
rect 6598 5468 6662 5472
rect 6598 5412 6602 5468
rect 6602 5412 6658 5468
rect 6658 5412 6662 5468
rect 6598 5408 6662 5412
rect 6678 5468 6742 5472
rect 6678 5412 6682 5468
rect 6682 5412 6738 5468
rect 6738 5412 6742 5468
rect 6678 5408 6742 5412
rect 1641 4924 1705 4928
rect 1641 4868 1645 4924
rect 1645 4868 1701 4924
rect 1701 4868 1705 4924
rect 1641 4864 1705 4868
rect 1721 4924 1785 4928
rect 1721 4868 1725 4924
rect 1725 4868 1781 4924
rect 1781 4868 1785 4924
rect 1721 4864 1785 4868
rect 1801 4924 1865 4928
rect 1801 4868 1805 4924
rect 1805 4868 1861 4924
rect 1861 4868 1865 4924
rect 1801 4864 1865 4868
rect 1881 4924 1945 4928
rect 1881 4868 1885 4924
rect 1885 4868 1941 4924
rect 1941 4868 1945 4924
rect 1881 4864 1945 4868
rect 3020 4924 3084 4928
rect 3020 4868 3024 4924
rect 3024 4868 3080 4924
rect 3080 4868 3084 4924
rect 3020 4864 3084 4868
rect 3100 4924 3164 4928
rect 3100 4868 3104 4924
rect 3104 4868 3160 4924
rect 3160 4868 3164 4924
rect 3100 4864 3164 4868
rect 3180 4924 3244 4928
rect 3180 4868 3184 4924
rect 3184 4868 3240 4924
rect 3240 4868 3244 4924
rect 3180 4864 3244 4868
rect 3260 4924 3324 4928
rect 3260 4868 3264 4924
rect 3264 4868 3320 4924
rect 3320 4868 3324 4924
rect 3260 4864 3324 4868
rect 4399 4924 4463 4928
rect 4399 4868 4403 4924
rect 4403 4868 4459 4924
rect 4459 4868 4463 4924
rect 4399 4864 4463 4868
rect 4479 4924 4543 4928
rect 4479 4868 4483 4924
rect 4483 4868 4539 4924
rect 4539 4868 4543 4924
rect 4479 4864 4543 4868
rect 4559 4924 4623 4928
rect 4559 4868 4563 4924
rect 4563 4868 4619 4924
rect 4619 4868 4623 4924
rect 4559 4864 4623 4868
rect 4639 4924 4703 4928
rect 4639 4868 4643 4924
rect 4643 4868 4699 4924
rect 4699 4868 4703 4924
rect 4639 4864 4703 4868
rect 5778 4924 5842 4928
rect 5778 4868 5782 4924
rect 5782 4868 5838 4924
rect 5838 4868 5842 4924
rect 5778 4864 5842 4868
rect 5858 4924 5922 4928
rect 5858 4868 5862 4924
rect 5862 4868 5918 4924
rect 5918 4868 5922 4924
rect 5858 4864 5922 4868
rect 5938 4924 6002 4928
rect 5938 4868 5942 4924
rect 5942 4868 5998 4924
rect 5998 4868 6002 4924
rect 5938 4864 6002 4868
rect 6018 4924 6082 4928
rect 6018 4868 6022 4924
rect 6022 4868 6078 4924
rect 6078 4868 6082 4924
rect 6018 4864 6082 4868
rect 2301 4380 2365 4384
rect 2301 4324 2305 4380
rect 2305 4324 2361 4380
rect 2361 4324 2365 4380
rect 2301 4320 2365 4324
rect 2381 4380 2445 4384
rect 2381 4324 2385 4380
rect 2385 4324 2441 4380
rect 2441 4324 2445 4380
rect 2381 4320 2445 4324
rect 2461 4380 2525 4384
rect 2461 4324 2465 4380
rect 2465 4324 2521 4380
rect 2521 4324 2525 4380
rect 2461 4320 2525 4324
rect 2541 4380 2605 4384
rect 2541 4324 2545 4380
rect 2545 4324 2601 4380
rect 2601 4324 2605 4380
rect 2541 4320 2605 4324
rect 3680 4380 3744 4384
rect 3680 4324 3684 4380
rect 3684 4324 3740 4380
rect 3740 4324 3744 4380
rect 3680 4320 3744 4324
rect 3760 4380 3824 4384
rect 3760 4324 3764 4380
rect 3764 4324 3820 4380
rect 3820 4324 3824 4380
rect 3760 4320 3824 4324
rect 3840 4380 3904 4384
rect 3840 4324 3844 4380
rect 3844 4324 3900 4380
rect 3900 4324 3904 4380
rect 3840 4320 3904 4324
rect 3920 4380 3984 4384
rect 3920 4324 3924 4380
rect 3924 4324 3980 4380
rect 3980 4324 3984 4380
rect 3920 4320 3984 4324
rect 5059 4380 5123 4384
rect 5059 4324 5063 4380
rect 5063 4324 5119 4380
rect 5119 4324 5123 4380
rect 5059 4320 5123 4324
rect 5139 4380 5203 4384
rect 5139 4324 5143 4380
rect 5143 4324 5199 4380
rect 5199 4324 5203 4380
rect 5139 4320 5203 4324
rect 5219 4380 5283 4384
rect 5219 4324 5223 4380
rect 5223 4324 5279 4380
rect 5279 4324 5283 4380
rect 5219 4320 5283 4324
rect 5299 4380 5363 4384
rect 5299 4324 5303 4380
rect 5303 4324 5359 4380
rect 5359 4324 5363 4380
rect 5299 4320 5363 4324
rect 6438 4380 6502 4384
rect 6438 4324 6442 4380
rect 6442 4324 6498 4380
rect 6498 4324 6502 4380
rect 6438 4320 6502 4324
rect 6518 4380 6582 4384
rect 6518 4324 6522 4380
rect 6522 4324 6578 4380
rect 6578 4324 6582 4380
rect 6518 4320 6582 4324
rect 6598 4380 6662 4384
rect 6598 4324 6602 4380
rect 6602 4324 6658 4380
rect 6658 4324 6662 4380
rect 6598 4320 6662 4324
rect 6678 4380 6742 4384
rect 6678 4324 6682 4380
rect 6682 4324 6738 4380
rect 6738 4324 6742 4380
rect 6678 4320 6742 4324
rect 1641 3836 1705 3840
rect 1641 3780 1645 3836
rect 1645 3780 1701 3836
rect 1701 3780 1705 3836
rect 1641 3776 1705 3780
rect 1721 3836 1785 3840
rect 1721 3780 1725 3836
rect 1725 3780 1781 3836
rect 1781 3780 1785 3836
rect 1721 3776 1785 3780
rect 1801 3836 1865 3840
rect 1801 3780 1805 3836
rect 1805 3780 1861 3836
rect 1861 3780 1865 3836
rect 1801 3776 1865 3780
rect 1881 3836 1945 3840
rect 1881 3780 1885 3836
rect 1885 3780 1941 3836
rect 1941 3780 1945 3836
rect 1881 3776 1945 3780
rect 3020 3836 3084 3840
rect 3020 3780 3024 3836
rect 3024 3780 3080 3836
rect 3080 3780 3084 3836
rect 3020 3776 3084 3780
rect 3100 3836 3164 3840
rect 3100 3780 3104 3836
rect 3104 3780 3160 3836
rect 3160 3780 3164 3836
rect 3100 3776 3164 3780
rect 3180 3836 3244 3840
rect 3180 3780 3184 3836
rect 3184 3780 3240 3836
rect 3240 3780 3244 3836
rect 3180 3776 3244 3780
rect 3260 3836 3324 3840
rect 3260 3780 3264 3836
rect 3264 3780 3320 3836
rect 3320 3780 3324 3836
rect 3260 3776 3324 3780
rect 4399 3836 4463 3840
rect 4399 3780 4403 3836
rect 4403 3780 4459 3836
rect 4459 3780 4463 3836
rect 4399 3776 4463 3780
rect 4479 3836 4543 3840
rect 4479 3780 4483 3836
rect 4483 3780 4539 3836
rect 4539 3780 4543 3836
rect 4479 3776 4543 3780
rect 4559 3836 4623 3840
rect 4559 3780 4563 3836
rect 4563 3780 4619 3836
rect 4619 3780 4623 3836
rect 4559 3776 4623 3780
rect 4639 3836 4703 3840
rect 4639 3780 4643 3836
rect 4643 3780 4699 3836
rect 4699 3780 4703 3836
rect 4639 3776 4703 3780
rect 5778 3836 5842 3840
rect 5778 3780 5782 3836
rect 5782 3780 5838 3836
rect 5838 3780 5842 3836
rect 5778 3776 5842 3780
rect 5858 3836 5922 3840
rect 5858 3780 5862 3836
rect 5862 3780 5918 3836
rect 5918 3780 5922 3836
rect 5858 3776 5922 3780
rect 5938 3836 6002 3840
rect 5938 3780 5942 3836
rect 5942 3780 5998 3836
rect 5998 3780 6002 3836
rect 5938 3776 6002 3780
rect 6018 3836 6082 3840
rect 6018 3780 6022 3836
rect 6022 3780 6078 3836
rect 6078 3780 6082 3836
rect 6018 3776 6082 3780
rect 2301 3292 2365 3296
rect 2301 3236 2305 3292
rect 2305 3236 2361 3292
rect 2361 3236 2365 3292
rect 2301 3232 2365 3236
rect 2381 3292 2445 3296
rect 2381 3236 2385 3292
rect 2385 3236 2441 3292
rect 2441 3236 2445 3292
rect 2381 3232 2445 3236
rect 2461 3292 2525 3296
rect 2461 3236 2465 3292
rect 2465 3236 2521 3292
rect 2521 3236 2525 3292
rect 2461 3232 2525 3236
rect 2541 3292 2605 3296
rect 2541 3236 2545 3292
rect 2545 3236 2601 3292
rect 2601 3236 2605 3292
rect 2541 3232 2605 3236
rect 3680 3292 3744 3296
rect 3680 3236 3684 3292
rect 3684 3236 3740 3292
rect 3740 3236 3744 3292
rect 3680 3232 3744 3236
rect 3760 3292 3824 3296
rect 3760 3236 3764 3292
rect 3764 3236 3820 3292
rect 3820 3236 3824 3292
rect 3760 3232 3824 3236
rect 3840 3292 3904 3296
rect 3840 3236 3844 3292
rect 3844 3236 3900 3292
rect 3900 3236 3904 3292
rect 3840 3232 3904 3236
rect 3920 3292 3984 3296
rect 3920 3236 3924 3292
rect 3924 3236 3980 3292
rect 3980 3236 3984 3292
rect 3920 3232 3984 3236
rect 5059 3292 5123 3296
rect 5059 3236 5063 3292
rect 5063 3236 5119 3292
rect 5119 3236 5123 3292
rect 5059 3232 5123 3236
rect 5139 3292 5203 3296
rect 5139 3236 5143 3292
rect 5143 3236 5199 3292
rect 5199 3236 5203 3292
rect 5139 3232 5203 3236
rect 5219 3292 5283 3296
rect 5219 3236 5223 3292
rect 5223 3236 5279 3292
rect 5279 3236 5283 3292
rect 5219 3232 5283 3236
rect 5299 3292 5363 3296
rect 5299 3236 5303 3292
rect 5303 3236 5359 3292
rect 5359 3236 5363 3292
rect 5299 3232 5363 3236
rect 6438 3292 6502 3296
rect 6438 3236 6442 3292
rect 6442 3236 6498 3292
rect 6498 3236 6502 3292
rect 6438 3232 6502 3236
rect 6518 3292 6582 3296
rect 6518 3236 6522 3292
rect 6522 3236 6578 3292
rect 6578 3236 6582 3292
rect 6518 3232 6582 3236
rect 6598 3292 6662 3296
rect 6598 3236 6602 3292
rect 6602 3236 6658 3292
rect 6658 3236 6662 3292
rect 6598 3232 6662 3236
rect 6678 3292 6742 3296
rect 6678 3236 6682 3292
rect 6682 3236 6738 3292
rect 6738 3236 6742 3292
rect 6678 3232 6742 3236
rect 1641 2748 1705 2752
rect 1641 2692 1645 2748
rect 1645 2692 1701 2748
rect 1701 2692 1705 2748
rect 1641 2688 1705 2692
rect 1721 2748 1785 2752
rect 1721 2692 1725 2748
rect 1725 2692 1781 2748
rect 1781 2692 1785 2748
rect 1721 2688 1785 2692
rect 1801 2748 1865 2752
rect 1801 2692 1805 2748
rect 1805 2692 1861 2748
rect 1861 2692 1865 2748
rect 1801 2688 1865 2692
rect 1881 2748 1945 2752
rect 1881 2692 1885 2748
rect 1885 2692 1941 2748
rect 1941 2692 1945 2748
rect 1881 2688 1945 2692
rect 3020 2748 3084 2752
rect 3020 2692 3024 2748
rect 3024 2692 3080 2748
rect 3080 2692 3084 2748
rect 3020 2688 3084 2692
rect 3100 2748 3164 2752
rect 3100 2692 3104 2748
rect 3104 2692 3160 2748
rect 3160 2692 3164 2748
rect 3100 2688 3164 2692
rect 3180 2748 3244 2752
rect 3180 2692 3184 2748
rect 3184 2692 3240 2748
rect 3240 2692 3244 2748
rect 3180 2688 3244 2692
rect 3260 2748 3324 2752
rect 3260 2692 3264 2748
rect 3264 2692 3320 2748
rect 3320 2692 3324 2748
rect 3260 2688 3324 2692
rect 4399 2748 4463 2752
rect 4399 2692 4403 2748
rect 4403 2692 4459 2748
rect 4459 2692 4463 2748
rect 4399 2688 4463 2692
rect 4479 2748 4543 2752
rect 4479 2692 4483 2748
rect 4483 2692 4539 2748
rect 4539 2692 4543 2748
rect 4479 2688 4543 2692
rect 4559 2748 4623 2752
rect 4559 2692 4563 2748
rect 4563 2692 4619 2748
rect 4619 2692 4623 2748
rect 4559 2688 4623 2692
rect 4639 2748 4703 2752
rect 4639 2692 4643 2748
rect 4643 2692 4699 2748
rect 4699 2692 4703 2748
rect 4639 2688 4703 2692
rect 5778 2748 5842 2752
rect 5778 2692 5782 2748
rect 5782 2692 5838 2748
rect 5838 2692 5842 2748
rect 5778 2688 5842 2692
rect 5858 2748 5922 2752
rect 5858 2692 5862 2748
rect 5862 2692 5918 2748
rect 5918 2692 5922 2748
rect 5858 2688 5922 2692
rect 5938 2748 6002 2752
rect 5938 2692 5942 2748
rect 5942 2692 5998 2748
rect 5998 2692 6002 2748
rect 5938 2688 6002 2692
rect 6018 2748 6082 2752
rect 6018 2692 6022 2748
rect 6022 2692 6078 2748
rect 6078 2692 6082 2748
rect 6018 2688 6082 2692
rect 2301 2204 2365 2208
rect 2301 2148 2305 2204
rect 2305 2148 2361 2204
rect 2361 2148 2365 2204
rect 2301 2144 2365 2148
rect 2381 2204 2445 2208
rect 2381 2148 2385 2204
rect 2385 2148 2441 2204
rect 2441 2148 2445 2204
rect 2381 2144 2445 2148
rect 2461 2204 2525 2208
rect 2461 2148 2465 2204
rect 2465 2148 2521 2204
rect 2521 2148 2525 2204
rect 2461 2144 2525 2148
rect 2541 2204 2605 2208
rect 2541 2148 2545 2204
rect 2545 2148 2601 2204
rect 2601 2148 2605 2204
rect 2541 2144 2605 2148
rect 3680 2204 3744 2208
rect 3680 2148 3684 2204
rect 3684 2148 3740 2204
rect 3740 2148 3744 2204
rect 3680 2144 3744 2148
rect 3760 2204 3824 2208
rect 3760 2148 3764 2204
rect 3764 2148 3820 2204
rect 3820 2148 3824 2204
rect 3760 2144 3824 2148
rect 3840 2204 3904 2208
rect 3840 2148 3844 2204
rect 3844 2148 3900 2204
rect 3900 2148 3904 2204
rect 3840 2144 3904 2148
rect 3920 2204 3984 2208
rect 3920 2148 3924 2204
rect 3924 2148 3980 2204
rect 3980 2148 3984 2204
rect 3920 2144 3984 2148
rect 5059 2204 5123 2208
rect 5059 2148 5063 2204
rect 5063 2148 5119 2204
rect 5119 2148 5123 2204
rect 5059 2144 5123 2148
rect 5139 2204 5203 2208
rect 5139 2148 5143 2204
rect 5143 2148 5199 2204
rect 5199 2148 5203 2204
rect 5139 2144 5203 2148
rect 5219 2204 5283 2208
rect 5219 2148 5223 2204
rect 5223 2148 5279 2204
rect 5279 2148 5283 2204
rect 5219 2144 5283 2148
rect 5299 2204 5363 2208
rect 5299 2148 5303 2204
rect 5303 2148 5359 2204
rect 5359 2148 5363 2204
rect 5299 2144 5363 2148
rect 6438 2204 6502 2208
rect 6438 2148 6442 2204
rect 6442 2148 6498 2204
rect 6498 2148 6502 2204
rect 6438 2144 6502 2148
rect 6518 2204 6582 2208
rect 6518 2148 6522 2204
rect 6522 2148 6578 2204
rect 6578 2148 6582 2204
rect 6518 2144 6582 2148
rect 6598 2204 6662 2208
rect 6598 2148 6602 2204
rect 6602 2148 6658 2204
rect 6658 2148 6662 2204
rect 6598 2144 6662 2148
rect 6678 2204 6742 2208
rect 6678 2148 6682 2204
rect 6682 2148 6738 2204
rect 6738 2148 6742 2204
rect 6678 2144 6742 2148
<< metal4 >>
rect 2293 7710 2613 7752
rect 1633 7104 1953 7664
rect 1633 7040 1641 7104
rect 1705 7050 1721 7104
rect 1785 7050 1801 7104
rect 1865 7050 1881 7104
rect 1945 7040 1953 7104
rect 1633 6814 1675 7040
rect 1911 6814 1953 7040
rect 1633 6016 1953 6814
rect 1633 5952 1641 6016
rect 1705 5952 1721 6016
rect 1785 5952 1801 6016
rect 1865 5952 1881 6016
rect 1945 5952 1953 6016
rect 1633 5691 1953 5952
rect 1633 5455 1675 5691
rect 1911 5455 1953 5691
rect 1633 4928 1953 5455
rect 1633 4864 1641 4928
rect 1705 4864 1721 4928
rect 1785 4864 1801 4928
rect 1865 4864 1881 4928
rect 1945 4864 1953 4928
rect 1633 4332 1953 4864
rect 1633 4096 1675 4332
rect 1911 4096 1953 4332
rect 1633 3840 1953 4096
rect 1633 3776 1641 3840
rect 1705 3776 1721 3840
rect 1785 3776 1801 3840
rect 1865 3776 1881 3840
rect 1945 3776 1953 3840
rect 1633 2973 1953 3776
rect 1633 2752 1675 2973
rect 1911 2752 1953 2973
rect 1633 2688 1641 2752
rect 1705 2688 1721 2737
rect 1785 2688 1801 2737
rect 1865 2688 1881 2737
rect 1945 2688 1953 2752
rect 1633 2128 1953 2688
rect 2293 7648 2335 7710
rect 2571 7648 2613 7710
rect 3672 7710 3992 7752
rect 2293 7584 2301 7648
rect 2605 7584 2613 7648
rect 2293 7474 2335 7584
rect 2571 7474 2613 7584
rect 2293 6560 2613 7474
rect 2293 6496 2301 6560
rect 2365 6496 2381 6560
rect 2445 6496 2461 6560
rect 2525 6496 2541 6560
rect 2605 6496 2613 6560
rect 2293 6351 2613 6496
rect 2293 6115 2335 6351
rect 2571 6115 2613 6351
rect 2293 5472 2613 6115
rect 2293 5408 2301 5472
rect 2365 5408 2381 5472
rect 2445 5408 2461 5472
rect 2525 5408 2541 5472
rect 2605 5408 2613 5472
rect 2293 4992 2613 5408
rect 2293 4756 2335 4992
rect 2571 4756 2613 4992
rect 2293 4384 2613 4756
rect 2293 4320 2301 4384
rect 2365 4320 2381 4384
rect 2445 4320 2461 4384
rect 2525 4320 2541 4384
rect 2605 4320 2613 4384
rect 2293 3633 2613 4320
rect 2293 3397 2335 3633
rect 2571 3397 2613 3633
rect 2293 3296 2613 3397
rect 2293 3232 2301 3296
rect 2365 3232 2381 3296
rect 2445 3232 2461 3296
rect 2525 3232 2541 3296
rect 2605 3232 2613 3296
rect 2293 2208 2613 3232
rect 2293 2144 2301 2208
rect 2365 2144 2381 2208
rect 2445 2144 2461 2208
rect 2525 2144 2541 2208
rect 2605 2144 2613 2208
rect 2293 2128 2613 2144
rect 3012 7104 3332 7664
rect 3012 7040 3020 7104
rect 3084 7050 3100 7104
rect 3164 7050 3180 7104
rect 3244 7050 3260 7104
rect 3324 7040 3332 7104
rect 3012 6814 3054 7040
rect 3290 6814 3332 7040
rect 3012 6016 3332 6814
rect 3012 5952 3020 6016
rect 3084 5952 3100 6016
rect 3164 5952 3180 6016
rect 3244 5952 3260 6016
rect 3324 5952 3332 6016
rect 3012 5691 3332 5952
rect 3012 5455 3054 5691
rect 3290 5455 3332 5691
rect 3012 4928 3332 5455
rect 3012 4864 3020 4928
rect 3084 4864 3100 4928
rect 3164 4864 3180 4928
rect 3244 4864 3260 4928
rect 3324 4864 3332 4928
rect 3012 4332 3332 4864
rect 3012 4096 3054 4332
rect 3290 4096 3332 4332
rect 3012 3840 3332 4096
rect 3012 3776 3020 3840
rect 3084 3776 3100 3840
rect 3164 3776 3180 3840
rect 3244 3776 3260 3840
rect 3324 3776 3332 3840
rect 3012 2973 3332 3776
rect 3012 2752 3054 2973
rect 3290 2752 3332 2973
rect 3012 2688 3020 2752
rect 3084 2688 3100 2737
rect 3164 2688 3180 2737
rect 3244 2688 3260 2737
rect 3324 2688 3332 2752
rect 3012 2128 3332 2688
rect 3672 7648 3714 7710
rect 3950 7648 3992 7710
rect 5051 7710 5371 7752
rect 3672 7584 3680 7648
rect 3984 7584 3992 7648
rect 3672 7474 3714 7584
rect 3950 7474 3992 7584
rect 3672 6560 3992 7474
rect 3672 6496 3680 6560
rect 3744 6496 3760 6560
rect 3824 6496 3840 6560
rect 3904 6496 3920 6560
rect 3984 6496 3992 6560
rect 3672 6351 3992 6496
rect 3672 6115 3714 6351
rect 3950 6115 3992 6351
rect 3672 5472 3992 6115
rect 3672 5408 3680 5472
rect 3744 5408 3760 5472
rect 3824 5408 3840 5472
rect 3904 5408 3920 5472
rect 3984 5408 3992 5472
rect 3672 4992 3992 5408
rect 3672 4756 3714 4992
rect 3950 4756 3992 4992
rect 3672 4384 3992 4756
rect 3672 4320 3680 4384
rect 3744 4320 3760 4384
rect 3824 4320 3840 4384
rect 3904 4320 3920 4384
rect 3984 4320 3992 4384
rect 3672 3633 3992 4320
rect 3672 3397 3714 3633
rect 3950 3397 3992 3633
rect 3672 3296 3992 3397
rect 3672 3232 3680 3296
rect 3744 3232 3760 3296
rect 3824 3232 3840 3296
rect 3904 3232 3920 3296
rect 3984 3232 3992 3296
rect 3672 2208 3992 3232
rect 3672 2144 3680 2208
rect 3744 2144 3760 2208
rect 3824 2144 3840 2208
rect 3904 2144 3920 2208
rect 3984 2144 3992 2208
rect 3672 2128 3992 2144
rect 4391 7104 4711 7664
rect 4391 7040 4399 7104
rect 4463 7050 4479 7104
rect 4543 7050 4559 7104
rect 4623 7050 4639 7104
rect 4703 7040 4711 7104
rect 4391 6814 4433 7040
rect 4669 6814 4711 7040
rect 4391 6016 4711 6814
rect 4391 5952 4399 6016
rect 4463 5952 4479 6016
rect 4543 5952 4559 6016
rect 4623 5952 4639 6016
rect 4703 5952 4711 6016
rect 4391 5691 4711 5952
rect 4391 5455 4433 5691
rect 4669 5455 4711 5691
rect 4391 4928 4711 5455
rect 4391 4864 4399 4928
rect 4463 4864 4479 4928
rect 4543 4864 4559 4928
rect 4623 4864 4639 4928
rect 4703 4864 4711 4928
rect 4391 4332 4711 4864
rect 4391 4096 4433 4332
rect 4669 4096 4711 4332
rect 4391 3840 4711 4096
rect 4391 3776 4399 3840
rect 4463 3776 4479 3840
rect 4543 3776 4559 3840
rect 4623 3776 4639 3840
rect 4703 3776 4711 3840
rect 4391 2973 4711 3776
rect 4391 2752 4433 2973
rect 4669 2752 4711 2973
rect 4391 2688 4399 2752
rect 4463 2688 4479 2737
rect 4543 2688 4559 2737
rect 4623 2688 4639 2737
rect 4703 2688 4711 2752
rect 4391 2128 4711 2688
rect 5051 7648 5093 7710
rect 5329 7648 5371 7710
rect 6430 7710 6750 7752
rect 5051 7584 5059 7648
rect 5363 7584 5371 7648
rect 5051 7474 5093 7584
rect 5329 7474 5371 7584
rect 5051 6560 5371 7474
rect 5051 6496 5059 6560
rect 5123 6496 5139 6560
rect 5203 6496 5219 6560
rect 5283 6496 5299 6560
rect 5363 6496 5371 6560
rect 5051 6351 5371 6496
rect 5051 6115 5093 6351
rect 5329 6115 5371 6351
rect 5051 5472 5371 6115
rect 5051 5408 5059 5472
rect 5123 5408 5139 5472
rect 5203 5408 5219 5472
rect 5283 5408 5299 5472
rect 5363 5408 5371 5472
rect 5051 4992 5371 5408
rect 5051 4756 5093 4992
rect 5329 4756 5371 4992
rect 5051 4384 5371 4756
rect 5051 4320 5059 4384
rect 5123 4320 5139 4384
rect 5203 4320 5219 4384
rect 5283 4320 5299 4384
rect 5363 4320 5371 4384
rect 5051 3633 5371 4320
rect 5051 3397 5093 3633
rect 5329 3397 5371 3633
rect 5051 3296 5371 3397
rect 5051 3232 5059 3296
rect 5123 3232 5139 3296
rect 5203 3232 5219 3296
rect 5283 3232 5299 3296
rect 5363 3232 5371 3296
rect 5051 2208 5371 3232
rect 5051 2144 5059 2208
rect 5123 2144 5139 2208
rect 5203 2144 5219 2208
rect 5283 2144 5299 2208
rect 5363 2144 5371 2208
rect 5051 2128 5371 2144
rect 5770 7104 6090 7664
rect 5770 7040 5778 7104
rect 5842 7050 5858 7104
rect 5922 7050 5938 7104
rect 6002 7050 6018 7104
rect 6082 7040 6090 7104
rect 5770 6814 5812 7040
rect 6048 6814 6090 7040
rect 5770 6016 6090 6814
rect 5770 5952 5778 6016
rect 5842 5952 5858 6016
rect 5922 5952 5938 6016
rect 6002 5952 6018 6016
rect 6082 5952 6090 6016
rect 5770 5691 6090 5952
rect 5770 5455 5812 5691
rect 6048 5455 6090 5691
rect 5770 4928 6090 5455
rect 5770 4864 5778 4928
rect 5842 4864 5858 4928
rect 5922 4864 5938 4928
rect 6002 4864 6018 4928
rect 6082 4864 6090 4928
rect 5770 4332 6090 4864
rect 5770 4096 5812 4332
rect 6048 4096 6090 4332
rect 5770 3840 6090 4096
rect 5770 3776 5778 3840
rect 5842 3776 5858 3840
rect 5922 3776 5938 3840
rect 6002 3776 6018 3840
rect 6082 3776 6090 3840
rect 5770 2973 6090 3776
rect 5770 2752 5812 2973
rect 6048 2752 6090 2973
rect 5770 2688 5778 2752
rect 5842 2688 5858 2737
rect 5922 2688 5938 2737
rect 6002 2688 6018 2737
rect 6082 2688 6090 2752
rect 5770 2128 6090 2688
rect 6430 7648 6472 7710
rect 6708 7648 6750 7710
rect 6430 7584 6438 7648
rect 6742 7584 6750 7648
rect 6430 7474 6472 7584
rect 6708 7474 6750 7584
rect 6430 6560 6750 7474
rect 6430 6496 6438 6560
rect 6502 6496 6518 6560
rect 6582 6496 6598 6560
rect 6662 6496 6678 6560
rect 6742 6496 6750 6560
rect 6430 6351 6750 6496
rect 6430 6115 6472 6351
rect 6708 6115 6750 6351
rect 6430 5472 6750 6115
rect 6867 5812 6933 5813
rect 6867 5748 6868 5812
rect 6932 5748 6933 5812
rect 6867 5747 6933 5748
rect 6870 5541 6930 5747
rect 6867 5540 6933 5541
rect 6867 5476 6868 5540
rect 6932 5476 6933 5540
rect 6867 5475 6933 5476
rect 6430 5408 6438 5472
rect 6502 5408 6518 5472
rect 6582 5408 6598 5472
rect 6662 5408 6678 5472
rect 6742 5408 6750 5472
rect 6430 4992 6750 5408
rect 6430 4756 6472 4992
rect 6708 4756 6750 4992
rect 6430 4384 6750 4756
rect 6430 4320 6438 4384
rect 6502 4320 6518 4384
rect 6582 4320 6598 4384
rect 6662 4320 6678 4384
rect 6742 4320 6750 4384
rect 6430 3633 6750 4320
rect 6430 3397 6472 3633
rect 6708 3397 6750 3633
rect 6430 3296 6750 3397
rect 6430 3232 6438 3296
rect 6502 3232 6518 3296
rect 6582 3232 6598 3296
rect 6662 3232 6678 3296
rect 6742 3232 6750 3296
rect 6430 2208 6750 3232
rect 6430 2144 6438 2208
rect 6502 2144 6518 2208
rect 6582 2144 6598 2208
rect 6662 2144 6678 2208
rect 6742 2144 6750 2208
rect 6430 2128 6750 2144
<< via4 >>
rect 1675 7040 1705 7050
rect 1705 7040 1721 7050
rect 1721 7040 1785 7050
rect 1785 7040 1801 7050
rect 1801 7040 1865 7050
rect 1865 7040 1881 7050
rect 1881 7040 1911 7050
rect 1675 6814 1911 7040
rect 1675 5455 1911 5691
rect 1675 4096 1911 4332
rect 1675 2752 1911 2973
rect 1675 2737 1705 2752
rect 1705 2737 1721 2752
rect 1721 2737 1785 2752
rect 1785 2737 1801 2752
rect 1801 2737 1865 2752
rect 1865 2737 1881 2752
rect 1881 2737 1911 2752
rect 2335 7648 2571 7710
rect 2335 7584 2365 7648
rect 2365 7584 2381 7648
rect 2381 7584 2445 7648
rect 2445 7584 2461 7648
rect 2461 7584 2525 7648
rect 2525 7584 2541 7648
rect 2541 7584 2571 7648
rect 2335 7474 2571 7584
rect 2335 6115 2571 6351
rect 2335 4756 2571 4992
rect 2335 3397 2571 3633
rect 3054 7040 3084 7050
rect 3084 7040 3100 7050
rect 3100 7040 3164 7050
rect 3164 7040 3180 7050
rect 3180 7040 3244 7050
rect 3244 7040 3260 7050
rect 3260 7040 3290 7050
rect 3054 6814 3290 7040
rect 3054 5455 3290 5691
rect 3054 4096 3290 4332
rect 3054 2752 3290 2973
rect 3054 2737 3084 2752
rect 3084 2737 3100 2752
rect 3100 2737 3164 2752
rect 3164 2737 3180 2752
rect 3180 2737 3244 2752
rect 3244 2737 3260 2752
rect 3260 2737 3290 2752
rect 3714 7648 3950 7710
rect 3714 7584 3744 7648
rect 3744 7584 3760 7648
rect 3760 7584 3824 7648
rect 3824 7584 3840 7648
rect 3840 7584 3904 7648
rect 3904 7584 3920 7648
rect 3920 7584 3950 7648
rect 3714 7474 3950 7584
rect 3714 6115 3950 6351
rect 3714 4756 3950 4992
rect 3714 3397 3950 3633
rect 4433 7040 4463 7050
rect 4463 7040 4479 7050
rect 4479 7040 4543 7050
rect 4543 7040 4559 7050
rect 4559 7040 4623 7050
rect 4623 7040 4639 7050
rect 4639 7040 4669 7050
rect 4433 6814 4669 7040
rect 4433 5455 4669 5691
rect 4433 4096 4669 4332
rect 4433 2752 4669 2973
rect 4433 2737 4463 2752
rect 4463 2737 4479 2752
rect 4479 2737 4543 2752
rect 4543 2737 4559 2752
rect 4559 2737 4623 2752
rect 4623 2737 4639 2752
rect 4639 2737 4669 2752
rect 5093 7648 5329 7710
rect 5093 7584 5123 7648
rect 5123 7584 5139 7648
rect 5139 7584 5203 7648
rect 5203 7584 5219 7648
rect 5219 7584 5283 7648
rect 5283 7584 5299 7648
rect 5299 7584 5329 7648
rect 5093 7474 5329 7584
rect 5093 6115 5329 6351
rect 5093 4756 5329 4992
rect 5093 3397 5329 3633
rect 5812 7040 5842 7050
rect 5842 7040 5858 7050
rect 5858 7040 5922 7050
rect 5922 7040 5938 7050
rect 5938 7040 6002 7050
rect 6002 7040 6018 7050
rect 6018 7040 6048 7050
rect 5812 6814 6048 7040
rect 5812 5455 6048 5691
rect 5812 4096 6048 4332
rect 5812 2752 6048 2973
rect 5812 2737 5842 2752
rect 5842 2737 5858 2752
rect 5858 2737 5922 2752
rect 5922 2737 5938 2752
rect 5938 2737 6002 2752
rect 6002 2737 6018 2752
rect 6018 2737 6048 2752
rect 6472 7648 6708 7710
rect 6472 7584 6502 7648
rect 6502 7584 6518 7648
rect 6518 7584 6582 7648
rect 6582 7584 6598 7648
rect 6598 7584 6662 7648
rect 6662 7584 6678 7648
rect 6678 7584 6708 7648
rect 6472 7474 6708 7584
rect 6472 6115 6708 6351
rect 6472 4756 6708 4992
rect 6472 3397 6708 3633
<< metal5 >>
rect 1056 7710 6750 7752
rect 1056 7474 2335 7710
rect 2571 7474 3714 7710
rect 3950 7474 5093 7710
rect 5329 7474 6472 7710
rect 6708 7474 6750 7710
rect 1056 7432 6750 7474
rect 1056 7050 6672 7092
rect 1056 6814 1675 7050
rect 1911 6814 3054 7050
rect 3290 6814 4433 7050
rect 4669 6814 5812 7050
rect 6048 6814 6672 7050
rect 1056 6772 6672 6814
rect 1056 6351 6750 6393
rect 1056 6115 2335 6351
rect 2571 6115 3714 6351
rect 3950 6115 5093 6351
rect 5329 6115 6472 6351
rect 6708 6115 6750 6351
rect 1056 6073 6750 6115
rect 1056 5691 6672 5733
rect 1056 5455 1675 5691
rect 1911 5455 3054 5691
rect 3290 5455 4433 5691
rect 4669 5455 5812 5691
rect 6048 5455 6672 5691
rect 1056 5413 6672 5455
rect 1056 4992 6750 5034
rect 1056 4756 2335 4992
rect 2571 4756 3714 4992
rect 3950 4756 5093 4992
rect 5329 4756 6472 4992
rect 6708 4756 6750 4992
rect 1056 4714 6750 4756
rect 1056 4332 6672 4374
rect 1056 4096 1675 4332
rect 1911 4096 3054 4332
rect 3290 4096 4433 4332
rect 4669 4096 5812 4332
rect 6048 4096 6672 4332
rect 1056 4054 6672 4096
rect 1056 3633 6750 3675
rect 1056 3397 2335 3633
rect 2571 3397 3714 3633
rect 3950 3397 5093 3633
rect 5329 3397 6472 3633
rect 6708 3397 6750 3633
rect 1056 3355 6750 3397
rect 1056 2973 6672 3015
rect 1056 2737 1675 2973
rect 1911 2737 3054 2973
rect 3290 2737 4433 2973
rect 4669 2737 5812 2973
rect 6048 2737 6672 2973
rect 1056 2695 6672 2737
use sky130_fd_sc_hd__or4_2  _09_
timestamp 0
transform 1 0 3036 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _10_
timestamp 0
transform -1 0 3220 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _11_
timestamp 0
transform 1 0 2392 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _12_
timestamp 0
transform 1 0 2852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _13_
timestamp 0
transform 1 0 2852 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _14_
timestamp 0
transform -1 0 4508 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _15_
timestamp 0
transform 1 0 4140 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _16_
timestamp 0
transform 1 0 4876 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _17_
timestamp 0
transform -1 0 5796 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _18_
timestamp 0
transform 1 0 5060 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _19_
timestamp 0
transform -1 0 2116 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _20_
timestamp 0
transform 1 0 2576 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _21_
timestamp 0
transform 1 0 2760 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _22_
timestamp 0
transform 1 0 4232 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _23_
timestamp 0
transform -1 0 4600 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _24_
timestamp 0
transform -1 0 4232 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _25_
timestamp 0
transform 1 0 2116 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3
timestamp 0
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_15
timestamp 0
transform 1 0 2484 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_21
timestamp 0
transform 1 0 3036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 0
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_29
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_35
timestamp 0
transform 1 0 4324 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 0
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 0
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 0
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_15
timestamp 0
transform 1 0 2484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_19
timestamp 0
transform 1 0 2852 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_23
timestamp 0
transform 1 0 3220 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_31
timestamp 0
transform 1 0 3956 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 0
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 0
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 0
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_3
timestamp 0
transform 1 0 1380 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_11
timestamp 0
transform 1 0 2116 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_26
timestamp 0
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_29
timestamp 0
transform 1 0 3772 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_37
timestamp 0
transform 1 0 4508 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_47
timestamp 0
transform 1 0 5428 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_51
timestamp 0
transform 1 0 5796 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_15
timestamp 0
transform 1 0 2484 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_22
timestamp 0
transform 1 0 3128 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_34
timestamp 0
transform 1 0 4232 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_46
timestamp 0
transform 1 0 5336 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_54
timestamp 0
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 0
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 0
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 0
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 0
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 0
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_53
timestamp 0
transform 1 0 5980 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 0
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 0
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 0
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_39
timestamp 0
transform 1 0 4692 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_50
timestamp 0
transform 1 0 5704 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_11
timestamp 0
transform 1 0 2116 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_17
timestamp 0
transform 1 0 2668 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_22
timestamp 0
transform 1 0 3128 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 0
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_53
timestamp 0
transform 1 0 5980 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_3
timestamp 0
transform 1 0 1380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_14
timestamp 0
transform 1 0 2392 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 0
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 0
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 0
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 0
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 0
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 0
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_29
timestamp 0
transform 1 0 3772 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_38
timestamp 0
transform 1 0 4600 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_50
timestamp 0
transform 1 0 5704 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_56
timestamp 0
transform 1 0 6256 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_9
timestamp 0
transform 1 0 1932 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_20
timestamp 0
transform 1 0 2944 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_27
timestamp 0
transform 1 0 3588 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_29
timestamp 0
transform 1 0 3772 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_37
timestamp 0
transform 1 0 4508 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_44
timestamp 0
transform 1 0 5152 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 0
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 0
transform 1 0 1656 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 0
transform -1 0 2944 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 0
transform -1 0 3588 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 0
transform -1 0 4876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 0
transform 1 0 3312 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 0
transform 1 0 6072 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 0
transform 1 0 6072 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 0
transform -1 0 1748 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 0
transform 1 0 1748 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output11
timestamp 0
transform 1 0 4600 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output12
timestamp 0
transform 1 0 3956 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 0
transform -1 0 3036 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 0
transform 1 0 3956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 0
transform 1 0 5980 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 0
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_10
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 0
transform -1 0 6624 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_11
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 0
transform -1 0 6624 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_12
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 0
transform -1 0 6624 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_13
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 0
transform -1 0 6624 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_14
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 0
transform -1 0 6624 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_15
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 0
transform -1 0 6624 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_16
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 0
transform -1 0 6624 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_17
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 0
transform -1 0 6624 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_18
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 0
transform -1 0 6624 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_19
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 0
transform -1 0 6624 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_20
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_21
timestamp 0
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_22
timestamp 0
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_23
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_24
timestamp 0
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_25
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_26
timestamp 0
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_27
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_28
timestamp 0
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_29
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_30
timestamp 0
transform 1 0 3680 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_31
timestamp 0
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
<< labels >>
rlabel metal1 s 3927 7616 3927 7616 4 VGND
rlabel metal1 s 3864 7072 3864 7072 4 VPWR
rlabel metal1 s 2622 3570 2622 3570 4 _00_
rlabel metal2 s 3174 3366 3174 3366 4 _01_
rlabel metal2 s 2806 3910 2806 3910 4 _02_
rlabel metal1 s 4692 3434 4692 3434 4 _03_
rlabel metal1 s 5106 3638 5106 3638 4 _04_
rlabel metal1 s 5566 3536 5566 3536 4 _05_
rlabel metal1 s 3726 6256 3726 6256 4 _06_
rlabel metal1 s 3220 5882 3220 5882 4 _07_
rlabel metal2 s 4646 6596 4646 6596 4 _08_
rlabel metal3 s 0 7488 800 7608 4 in[0]
port 3 nsew
rlabel metal3 s 1096 6868 1096 6868 4 in[1]
rlabel metal2 s 2714 8279 2714 8279 4 in[2]
rlabel metal2 s 3358 8279 3358 8279 4 in[3]
rlabel metal2 s 4554 1588 4554 1588 4 in[4]
rlabel metal2 s 3266 1588 3266 1588 4 in[5]
rlabel metal2 s 6302 4369 6302 4369 4 in[6]
rlabel metal2 s 6302 5729 6302 5729 4 in[7]
rlabel metal1 s 1610 6222 1610 6222 4 net1
rlabel metal1 s 1794 5712 1794 5712 4 net10
rlabel metal1 s 4692 6970 4692 6970 4 net11
rlabel metal1 s 4002 6426 4002 6426 4 net12
rlabel metal1 s 2944 2414 2944 2414 4 net13
rlabel metal1 s 3726 2414 3726 2414 4 net14
rlabel metal1 s 5888 3502 5888 3502 4 net15
rlabel metal1 s 5658 5168 5658 5168 4 net16
rlabel metal1 s 1978 6290 1978 6290 4 net2
rlabel metal1 s 2852 6290 2852 6290 4 net3
rlabel metal1 s 3680 6426 3680 6426 4 net4
rlabel metal1 s 2530 3468 2530 3468 4 net5
rlabel metal1 s 4140 3638 4140 3638 4 net6
rlabel metal1 s 4002 3536 4002 3536 4 net7
rlabel metal1 s 5382 5202 5382 5202 4 net8
rlabel metal1 s 1702 5644 1702 5644 4 net9
rlabel metal1 s 1380 5882 1380 5882 4 out[0]
rlabel metal3 s 1326 5508 1326 5508 4 out[1]
rlabel metal2 s 4830 8347 4830 8347 4 out[2]
rlabel metal1 s 4140 7514 4140 7514 4 out[3]
rlabel metal2 s 2622 959 2622 959 4 out[4]
rlabel metal2 s 3910 959 3910 959 4 out[5]
rlabel metal2 s 6210 3417 6210 3417 4 out[6]
rlabel metal1 s 6164 4998 6164 4998 4 out[7]
flabel metal5 s 1056 7432 6750 7752 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 6073 6750 6393 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 4714 6750 5034 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 3355 6750 3675 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal4 s 6430 2128 6750 7752 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 5051 2128 5371 7752 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 3672 2128 3992 7752 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 2293 2128 2613 7752 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal5 s 1056 6772 6672 7092 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 5413 6672 5733 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 4054 6672 4374 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 2695 6672 3015 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal4 s 5770 2128 6090 7664 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 4391 2128 4711 7664 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 3012 2128 3332 7664 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 1633 2128 1953 7664 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal3 s 400 7548 400 7548 0 FreeSans 600 0 0 0 in[0]
flabel metal3 s 0 6808 800 6928 0 FreeSans 600 0 0 0 in[1]
port 4 nsew
flabel metal2 s 2594 9077 2650 9877 0 FreeSans 280 90 0 0 in[2]
port 5 nsew
flabel metal2 s 3238 9077 3294 9877 0 FreeSans 280 90 0 0 in[3]
port 6 nsew
flabel metal2 s 4526 0 4582 800 0 FreeSans 280 90 0 0 in[4]
port 7 nsew
flabel metal2 s 3238 0 3294 800 0 FreeSans 280 90 0 0 in[5]
port 8 nsew
flabel metal3 s 6933 4088 7733 4208 0 FreeSans 600 0 0 0 in[6]
port 9 nsew
flabel metal3 s 6933 5448 7733 5568 0 FreeSans 600 0 0 0 in[7]
port 10 nsew
flabel metal3 s 0 6128 800 6248 0 FreeSans 600 0 0 0 out[0]
port 11 nsew
flabel metal3 s 0 5448 800 5568 0 FreeSans 600 0 0 0 out[1]
port 12 nsew
flabel metal2 s 4526 9077 4582 9877 0 FreeSans 280 90 0 0 out[2]
port 13 nsew
flabel metal2 s 3882 9077 3938 9877 0 FreeSans 280 90 0 0 out[3]
port 14 nsew
flabel metal2 s 2594 0 2650 800 0 FreeSans 280 90 0 0 out[4]
port 15 nsew
flabel metal2 s 3882 0 3938 800 0 FreeSans 280 90 0 0 out[5]
port 16 nsew
flabel metal3 s 6933 3408 7733 3528 0 FreeSans 600 0 0 0 out[6]
port 17 nsew
flabel metal3 s 6933 4768 7733 4888 0 FreeSans 600 0 0 0 out[7]
port 18 nsew
<< properties >>
string FIXED_BBOX 0 0 7733 9877
<< end >>
